* NGSPICE file created from CaravelHost.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

.subckt CaravelHost caravel_uart_rx caravel_uart_tx caravel_wb_ack_i caravel_wb_adr_o[0]
+ caravel_wb_adr_o[10] caravel_wb_adr_o[11] caravel_wb_adr_o[12] caravel_wb_adr_o[13]
+ caravel_wb_adr_o[14] caravel_wb_adr_o[15] caravel_wb_adr_o[16] caravel_wb_adr_o[17]
+ caravel_wb_adr_o[18] caravel_wb_adr_o[19] caravel_wb_adr_o[1] caravel_wb_adr_o[20]
+ caravel_wb_adr_o[21] caravel_wb_adr_o[22] caravel_wb_adr_o[23] caravel_wb_adr_o[24]
+ caravel_wb_adr_o[25] caravel_wb_adr_o[26] caravel_wb_adr_o[27] caravel_wb_adr_o[2]
+ caravel_wb_adr_o[3] caravel_wb_adr_o[4] caravel_wb_adr_o[5] caravel_wb_adr_o[6]
+ caravel_wb_adr_o[7] caravel_wb_adr_o[8] caravel_wb_adr_o[9] caravel_wb_cyc_o caravel_wb_data_i[0]
+ caravel_wb_data_i[10] caravel_wb_data_i[11] caravel_wb_data_i[12] caravel_wb_data_i[13]
+ caravel_wb_data_i[14] caravel_wb_data_i[15] caravel_wb_data_i[16] caravel_wb_data_i[17]
+ caravel_wb_data_i[18] caravel_wb_data_i[19] caravel_wb_data_i[1] caravel_wb_data_i[20]
+ caravel_wb_data_i[21] caravel_wb_data_i[22] caravel_wb_data_i[23] caravel_wb_data_i[24]
+ caravel_wb_data_i[25] caravel_wb_data_i[26] caravel_wb_data_i[27] caravel_wb_data_i[28]
+ caravel_wb_data_i[29] caravel_wb_data_i[2] caravel_wb_data_i[30] caravel_wb_data_i[31]
+ caravel_wb_data_i[3] caravel_wb_data_i[4] caravel_wb_data_i[5] caravel_wb_data_i[6]
+ caravel_wb_data_i[7] caravel_wb_data_i[8] caravel_wb_data_i[9] caravel_wb_data_o[0]
+ caravel_wb_data_o[10] caravel_wb_data_o[11] caravel_wb_data_o[12] caravel_wb_data_o[13]
+ caravel_wb_data_o[14] caravel_wb_data_o[15] caravel_wb_data_o[16] caravel_wb_data_o[17]
+ caravel_wb_data_o[18] caravel_wb_data_o[19] caravel_wb_data_o[1] caravel_wb_data_o[20]
+ caravel_wb_data_o[21] caravel_wb_data_o[22] caravel_wb_data_o[23] caravel_wb_data_o[24]
+ caravel_wb_data_o[25] caravel_wb_data_o[26] caravel_wb_data_o[27] caravel_wb_data_o[28]
+ caravel_wb_data_o[29] caravel_wb_data_o[2] caravel_wb_data_o[30] caravel_wb_data_o[31]
+ caravel_wb_data_o[3] caravel_wb_data_o[4] caravel_wb_data_o[5] caravel_wb_data_o[6]
+ caravel_wb_data_o[7] caravel_wb_data_o[8] caravel_wb_data_o[9] caravel_wb_error_i
+ caravel_wb_sel_o[0] caravel_wb_sel_o[1] caravel_wb_sel_o[2] caravel_wb_sel_o[3]
+ caravel_wb_stall_i caravel_wb_stb_o caravel_wb_we_o core0Index[0] core0Index[1]
+ core0Index[2] core0Index[3] core0Index[4] core0Index[5] core0Index[6] core0Index[7]
+ core1Index[0] core1Index[1] core1Index[2] core1Index[3] core1Index[4] core1Index[5]
+ core1Index[6] core1Index[7] manufacturerID[0] manufacturerID[10] manufacturerID[1]
+ manufacturerID[2] manufacturerID[3] manufacturerID[4] manufacturerID[5] manufacturerID[6]
+ manufacturerID[7] manufacturerID[8] manufacturerID[9] partID[0] partID[10] partID[11]
+ partID[12] partID[13] partID[14] partID[15] partID[1] partID[2] partID[3] partID[4]
+ partID[5] partID[6] partID[7] partID[8] partID[9] vccd1 versionID[0] versionID[1]
+ versionID[2] versionID[3] vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_data_i[0] wbs_data_i[10] wbs_data_i[11] wbs_data_i[12] wbs_data_i[13] wbs_data_i[14]
+ wbs_data_i[15] wbs_data_i[16] wbs_data_i[17] wbs_data_i[18] wbs_data_i[19] wbs_data_i[1]
+ wbs_data_i[20] wbs_data_i[21] wbs_data_i[22] wbs_data_i[23] wbs_data_i[24] wbs_data_i[25]
+ wbs_data_i[26] wbs_data_i[27] wbs_data_i[28] wbs_data_i[29] wbs_data_i[2] wbs_data_i[30]
+ wbs_data_i[31] wbs_data_i[3] wbs_data_i[4] wbs_data_i[5] wbs_data_i[6] wbs_data_i[7]
+ wbs_data_i[8] wbs_data_i[9] wbs_data_o[0] wbs_data_o[10] wbs_data_o[11] wbs_data_o[12]
+ wbs_data_o[13] wbs_data_o[14] wbs_data_o[15] wbs_data_o[16] wbs_data_o[17] wbs_data_o[18]
+ wbs_data_o[19] wbs_data_o[1] wbs_data_o[20] wbs_data_o[21] wbs_data_o[22] wbs_data_o[23]
+ wbs_data_o[24] wbs_data_o[25] wbs_data_o[26] wbs_data_o[27] wbs_data_o[28] wbs_data_o[29]
+ wbs_data_o[2] wbs_data_o[30] wbs_data_o[31] wbs_data_o[3] wbs_data_o[4] wbs_data_o[5]
+ wbs_data_o[6] wbs_data_o[7] wbs_data_o[8] wbs_data_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6914_ _6914_/A vssd1 vssd1 vccd1 vccd1 _7669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6845_ _6849_/B _6845_/B _6859_/C vssd1 vssd1 vccd1 vccd1 _6846_/A sky130_fd_sc_hd__and3b_1
XFILLER_23_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3988_ _3644_/X _7523_/Q _3994_/S vssd1 vssd1 vccd1 vccd1 _3989_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6776_ _6100_/Y _6101_/X _6775_/X _6157_/C _6164_/C vssd1 vssd1 vccd1 vccd1 _6779_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_23_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4609_ _4609_/A vssd1 vssd1 vccd1 vccd1 _7257_/D sky130_fd_sc_hd__clkbuf_1
X_5589_ _7080_/Q _5588_/X _5380_/C _5587_/B vssd1 vssd1 vccd1 vccd1 _5590_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7328_ _7525_/CLK _7328_/D vssd1 vssd1 vccd1 vccd1 _7328_/Q sky130_fd_sc_hd__dfxtp_4
X_7259_ _7259_/CLK _7259_/D vssd1 vssd1 vccd1 vccd1 _7259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3084_ clkbuf_0__3084_/X vssd1 vssd1 vccd1 vccd1 _6301__439/A sky130_fd_sc_hd__clkbuf_16
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6940__30 _6941__31/A vssd1 vssd1 vccd1 vccd1 _7686_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _5555_/A _4966_/B vssd1 vssd1 vccd1 vccd1 _4961_/A sky130_fd_sc_hd__and2_1
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3911_ _3911_/A vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__clkbuf_4
X_4891_ _4891_/A vssd1 vssd1 vccd1 vccd1 _7076_/D sky130_fd_sc_hd__clkbuf_1
X_3842_ _4121_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _3858_/S sky130_fd_sc_hd__or2_4
X_6561_ _6561_/A vssd1 vssd1 vccd1 vccd1 _6589_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3773_ _3773_/A vssd1 vssd1 vccd1 vccd1 _7607_/D sky130_fd_sc_hd__clkbuf_1
X_5512_ _7034_/A vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6492_ _7508_/Q _6492_/B _6492_/C vssd1 vssd1 vccd1 vccd1 _6505_/B sky130_fd_sc_hd__and3_1
X_5443_ _5493_/S input33/X _5449_/A _6481_/A vssd1 vssd1 vccd1 vccd1 _5443_/X sky130_fd_sc_hd__a22o_1
X_5374_ _5374_/A vssd1 vssd1 vccd1 vccd1 _5374_/X sky130_fd_sc_hd__clkbuf_1
X_7113_ _7113_/CLK _7113_/D vssd1 vssd1 vccd1 vccd1 _7113_/Q sky130_fd_sc_hd__dfxtp_1
X_4325_ _7327_/Q vssd1 vssd1 vccd1 vccd1 _4325_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4256_ _4255_/X _7394_/Q _4262_/S vssd1 vssd1 vccd1 vccd1 _4257_/A sky130_fd_sc_hd__mux2_1
X_7044_ _5496_/A _7044_/D vssd1 vssd1 vccd1 vccd1 _7044_/Q sky130_fd_sc_hd__dfxtp_1
X_4187_ _4112_/X _7418_/Q _4191_/S vssd1 vssd1 vccd1 vccd1 _4188_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2956_ _6037_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2956_/X sky130_fd_sc_hd__clkbuf_16
X_6828_ _6828_/A vssd1 vssd1 vccd1 vccd1 _7644_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6400__519 _6400__519/A vssd1 vssd1 vccd1 vccd1 _7461_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6292__432 _6292__432/A vssd1 vssd1 vccd1 vccd1 _7374_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2722_ clkbuf_0__2722_/X vssd1 vssd1 vccd1 vccd1 _5736__284/A sky130_fd_sc_hd__clkbuf_16
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6301__439 _6301__439/A vssd1 vssd1 vccd1 vccd1 _7381_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__3281_ clkbuf_0__3281_/X vssd1 vssd1 vccd1 vccd1 _6700__139/A sky130_fd_sc_hd__clkbuf_16
XFILLER_52_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5090_ _7198_/Q _5090_/B vssd1 vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__and2_1
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4110_ _4109_/X _7451_/Q _4110_/S vssd1 vssd1 vccd1 vccd1 _4111_/A sky130_fd_sc_hd__mux2_1
X_4041_ _4056_/S vssd1 vssd1 vccd1 vccd1 _4050_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5992_ _7224_/Q _5814_/A _5990_/X _5991_/X vssd1 vssd1 vccd1 vccd1 _7224_/D sky130_fd_sc_hd__o211a_1
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _4943_/A vssd1 vssd1 vccd1 vccd1 _7041_/D sky130_fd_sc_hd__clkbuf_1
X_7731_ _7731_/CLK _7731_/D vssd1 vssd1 vccd1 vccd1 _7731_/Q sky130_fd_sc_hd__dfxtp_1
X_7662_ _7727_/CLK _7662_/D vssd1 vssd1 vccd1 vccd1 _7662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4874_ _4834_/X _7109_/Q _4874_/S vssd1 vssd1 vccd1 vccd1 _4875_/A sky130_fd_sc_hd__mux2_1
X_6613_ _7516_/Q _7497_/Q _6525_/A _6610_/Y _6515_/B vssd1 vssd1 vccd1 vccd1 _6615_/B
+ sky130_fd_sc_hd__a2111o_1
X_7593_ _7593_/CLK _7593_/D vssd1 vssd1 vccd1 vccd1 _7593_/Q sky130_fd_sc_hd__dfxtp_1
X_3825_ _3840_/S vssd1 vssd1 vccd1 vccd1 _3834_/S sky130_fd_sc_hd__clkbuf_4
X_6762__14 _6762__14/A vssd1 vssd1 vccd1 vccd1 _7633_/CLK sky130_fd_sc_hd__inv_2
X_3756_ _3756_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _4361_/B sky130_fd_sc_hd__nand2_1
X_6544_ _6553_/C _6583_/C _6544_/C vssd1 vssd1 vccd1 vccd1 _6544_/X sky130_fd_sc_hd__and3b_1
XFILLER_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6475_ _6469_/X _6470_/Y _6473_/Y _6474_/X vssd1 vssd1 vccd1 vccd1 _6475_/X sky130_fd_sc_hd__a211o_1
XFILLER_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3687_ _3687_/A vssd1 vssd1 vccd1 vccd1 _7676_/D sky130_fd_sc_hd__clkbuf_1
X_5426_ _5422_/X _5424_/X _5425_/X _5415_/A _5205_/A vssd1 vssd1 vccd1 vccd1 _5433_/B
+ sky130_fd_sc_hd__o221a_1
X_6356__484 _6356__484/A vssd1 vssd1 vccd1 vccd1 _7426_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5357_ _7119_/Q _7167_/Q _5421_/S vssd1 vssd1 vccd1 vccd1 _5358_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_4 _3603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5288_ _7529_/Q _7109_/Q _7561_/Q _7125_/Q _5173_/A _5171_/X vssd1 vssd1 vccd1 vccd1
+ _5289_/B sky130_fd_sc_hd__mux4_1
X_4308_ _4220_/X _7373_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4309_/A sky130_fd_sc_hd__mux2_1
X_4239_ _4239_/A _4642_/B vssd1 vssd1 vccd1 vccd1 _4262_/S sky130_fd_sc_hd__or2_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7027_ _6913_/A _6119_/B _7033_/S vssd1 vssd1 vccd1 vccd1 _7028_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3086_ _6308_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3086_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6755__8 _6756__9/A vssd1 vssd1 vccd1 vccd1 _7627_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2636_ clkbuf_0__2636_/X vssd1 vssd1 vccd1 vccd1 _5522__193/A sky130_fd_sc_hd__clkbuf_16
XFILLER_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4590_ _4238_/X _7265_/Q _4598_/S vssd1 vssd1 vccd1 vccd1 _4591_/A sky130_fd_sc_hd__mux2_1
X_3610_ _3610_/A vssd1 vssd1 vccd1 vccd1 _6915_/A sky130_fd_sc_hd__clkbuf_16
X_3541_ _7668_/Q vssd1 vssd1 vccd1 vccd1 _3920_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6260_ _6260_/A vssd1 vssd1 vccd1 vccd1 _6260_/X sky130_fd_sc_hd__buf_1
X_3472_ _7318_/Q vssd1 vssd1 vccd1 vccd1 _4095_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5804__294 _5804__294/A vssd1 vssd1 vccd1 vccd1 _7212_/CLK sky130_fd_sc_hd__inv_2
X_5211_ _5270_/A vssd1 vssd1 vccd1 vccd1 _5362_/S sky130_fd_sc_hd__clkbuf_4
X_5142_ _5262_/A vssd1 vssd1 vccd1 vccd1 _5356_/A sky130_fd_sc_hd__buf_2
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5073_ _5073_/A _5079_/B vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__and2_1
X_4024_ _4024_/A vssd1 vssd1 vccd1 vccd1 _7487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5975_ _5973_/X _5974_/X _5995_/S vssd1 vssd1 vccd1 vccd1 _5975_/X sky130_fd_sc_hd__mux2_2
XFILLER_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7714_ _7714_/CLK _7714_/D vssd1 vssd1 vccd1 vccd1 _7714_/Q sky130_fd_sc_hd__dfxtp_1
X_4926_ _7049_/Q _4572_/A _4928_/S vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__2724_ _5738_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2724_/X sky130_fd_sc_hd__clkbuf_16
X_4857_ _4857_/A vssd1 vssd1 vccd1 vccd1 _7117_/D sky130_fd_sc_hd__clkbuf_1
X_7645_ _7652_/CLK _7645_/D vssd1 vssd1 vccd1 vccd1 _7645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7576_ _7576_/CLK _7576_/D vssd1 vssd1 vccd1 vccd1 _7576_/Q sky130_fd_sc_hd__dfxtp_1
X_3808_ _7594_/Q _3807_/X _3811_/S vssd1 vssd1 vccd1 vccd1 _3809_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6527_ _6532_/C _6566_/A _6526_/X _5991_/X vssd1 vssd1 vccd1 vccd1 _7498_/D sky130_fd_sc_hd__o211a_1
X_4788_ _7144_/Q _4566_/A _4794_/S vssd1 vssd1 vccd1 vccd1 _4789_/A sky130_fd_sc_hd__mux2_1
X_3739_ _3738_/X _7619_/Q _3745_/S vssd1 vssd1 vccd1 vccd1 _3740_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6458_ _6463_/A _6458_/B vssd1 vssd1 vccd1 vccd1 _6459_/B sky130_fd_sc_hd__xnor2_1
X_6389_ _6395_/A vssd1 vssd1 vccd1 vccd1 _6389_/X sky130_fd_sc_hd__buf_1
XFILLER_0_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5409_ _5381_/Y _5394_/X _5407_/X _5441_/D _6133_/A vssd1 vssd1 vccd1 vccd1 _5410_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_102_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6040__322 _6042__324/A vssd1 vssd1 vccd1 vccd1 _7248_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5760_ _5004_/A _7191_/Q _5764_/S vssd1 vssd1 vccd1 vccd1 _5761_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4711_ _4711_/A vssd1 vssd1 vccd1 vccd1 _7179_/D sky130_fd_sc_hd__clkbuf_1
X_4642_ _4642_/A _4642_/B vssd1 vssd1 vccd1 vccd1 _4658_/S sky130_fd_sc_hd__or2_2
X_7430_ _7430_/CLK _7430_/D vssd1 vssd1 vccd1 vccd1 _7430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ _4572_/X _7270_/Q _4576_/S vssd1 vssd1 vccd1 vccd1 _4574_/A sky130_fd_sc_hd__mux2_1
X_7361_ _7361_/CLK _7361_/D vssd1 vssd1 vccd1 vccd1 _7361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3524_ _3524_/A vssd1 vssd1 vccd1 vccd1 _7713_/D sky130_fd_sc_hd__clkbuf_1
X_7292_ _7292_/CLK _7292_/D vssd1 vssd1 vccd1 vccd1 _7292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5125_ _7096_/Q _7097_/Q _5645_/B _5125_/D vssd1 vssd1 vccd1 vccd1 _5126_/D sky130_fd_sc_hd__or4_1
X_5056_ _5056_/A vssd1 vssd1 vccd1 vccd1 _5056_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4007_ _7494_/Q _3585_/X _4013_/S vssd1 vssd1 vccd1 vccd1 _4008_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5958_ _7215_/Q _7041_/Q _7263_/Q _7255_/Q _5841_/X _5913_/X vssd1 vssd1 vccd1 vccd1
+ _5958_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4909_ _4909_/A vssd1 vssd1 vccd1 vccd1 _7057_/D sky130_fd_sc_hd__clkbuf_1
X_5889_ _7624_/Q _7616_/Q _7600_/Q _7592_/Q _4484_/X _4477_/A vssd1 vssd1 vccd1 vccd1
+ _5890_/B sky130_fd_sc_hd__mux4_2
Xclkbuf_0__2707_ _5651_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2707_/X sky130_fd_sc_hd__clkbuf_16
X_7628_ _7628_/CLK _7628_/D vssd1 vssd1 vccd1 vccd1 _7628_/Q sky130_fd_sc_hd__dfxtp_1
X_7559_ _7559_/CLK _7559_/D vssd1 vssd1 vccd1 vccd1 _7559_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2638_ _5530_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2638_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6369__494 _6369__494/A vssd1 vssd1 vccd1 vccd1 _7436_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6947__36 _6948__37/A vssd1 vssd1 vccd1 vccd1 _7692_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3101_ clkbuf_0__3101_/X vssd1 vssd1 vccd1 vccd1 _6395_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_113_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6861_ _6889_/B _6878_/D vssd1 vssd1 vccd1 vccd1 _6876_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6047__328 _6048__329/A vssd1 vssd1 vccd1 vccd1 _7254_/CLK sky130_fd_sc_hd__inv_2
X_5812_ _6236_/C _6607_/B vssd1 vssd1 vccd1 vccd1 _5833_/A sky130_fd_sc_hd__and2_2
XFILLER_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6792_ _6792_/A _6792_/B _6792_/C _6792_/D vssd1 vssd1 vccd1 vccd1 _6792_/Y sky130_fd_sc_hd__nand4_1
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4625_ _4640_/S vssd1 vssd1 vccd1 vccd1 _4634_/S sky130_fd_sc_hd__buf_2
X_7413_ _7413_/CLK _7413_/D vssd1 vssd1 vccd1 vccd1 _7413_/Q sky130_fd_sc_hd__dfxtp_1
X_4556_ _7278_/Q _3920_/A _4558_/S vssd1 vssd1 vccd1 vccd1 _4557_/A sky130_fd_sc_hd__mux2_1
X_7344_ _7344_/CLK _7344_/D vssd1 vssd1 vccd1 vccd1 _7344_/Q sky130_fd_sc_hd__dfxtp_1
X_3507_ _7274_/Q vssd1 vssd1 vccd1 vccd1 _3510_/B sky130_fd_sc_hd__inv_2
XFILLER_116_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4487_ _4487_/A vssd1 vssd1 vccd1 vccd1 _7310_/D sky130_fd_sc_hd__clkbuf_1
X_7275_ _5496_/A _7275_/D vssd1 vssd1 vccd1 vccd1 _7275_/Q sky130_fd_sc_hd__dfxtp_1
X_6226_ _6226_/A vssd1 vssd1 vccd1 vccd1 _7325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6157_/A _6157_/B _6157_/C _6774_/A vssd1 vssd1 vccd1 vccd1 _6165_/C sky130_fd_sc_hd__or4_1
XFILLER_111_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _7044_/Q vssd1 vssd1 vccd1 vccd1 _5592_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_85_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6088_ _6908_/A _3513_/X _5535_/B vssd1 vssd1 vccd1 vccd1 _6797_/A sky130_fd_sc_hd__a21oi_2
X_5039_ _5039_/A vssd1 vssd1 vccd1 vccd1 _5039_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6731__164 _6731__164/A vssd1 vssd1 vccd1 vccd1 _7608_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__2953_ clkbuf_0__2953_/X vssd1 vssd1 vccd1 vccd1 _6031_/A sky130_fd_sc_hd__clkbuf_16
Xoutput97 _5076_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[13] sky130_fd_sc_hd__buf_2
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XCaravelHost_203 vssd1 vssd1 vccd1 vccd1 CaravelHost_203/HI core1Index[3] sky130_fd_sc_hd__conb_1
XFILLER_117_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_225 vssd1 vssd1 vccd1 vccd1 CaravelHost_225/HI partID[13] sky130_fd_sc_hd__conb_1
XCaravelHost_236 vssd1 vssd1 vccd1 vccd1 partID[10] CaravelHost_236/LO sky130_fd_sc_hd__conb_1
XCaravelHost_214 vssd1 vssd1 vccd1 vccd1 CaravelHost_214/HI manufacturerID[6] sky130_fd_sc_hd__conb_1
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4410_ _7342_/Q _4334_/X _4410_/S vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__mux2_1
X_5390_ _7438_/Q _4396_/X _5389_/X vssd1 vssd1 vccd1 vccd1 _5390_/X sky130_fd_sc_hd__o21a_1
X_4341_ _7361_/Q _4340_/X _4344_/S vssd1 vssd1 vccd1 vccd1 _4342_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4272_ _4272_/A vssd1 vssd1 vccd1 vccd1 _7389_/D sky130_fd_sc_hd__clkbuf_1
X_7060_ _7060_/CLK _7060_/D vssd1 vssd1 vccd1 vccd1 _7060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6350__479 _6350__479/A vssd1 vssd1 vccd1 vccd1 _7421_/CLK sky130_fd_sc_hd__inv_2
X_6011_ _7225_/Q _5814_/A _6010_/X _5991_/X vssd1 vssd1 vccd1 vccd1 _7225_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5695__250 _5698__253/A vssd1 vssd1 vccd1 vccd1 _7144_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6913_ _6913_/A _6923_/B vssd1 vssd1 vccd1 vccd1 _6914_/A sky130_fd_sc_hd__and2_1
XFILLER_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6844_ _6847_/C _6843_/C _7648_/Q vssd1 vssd1 vccd1 vccd1 _6845_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6674__118 _6674__118/A vssd1 vssd1 vccd1 vccd1 _7562_/CLK sky130_fd_sc_hd__inv_2
X_3987_ _3987_/A vssd1 vssd1 vccd1 vccd1 _7524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6775_ _6775_/A _6775_/B vssd1 vssd1 vccd1 vccd1 _6775_/X sky130_fd_sc_hd__or2_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5657_ _5663_/A vssd1 vssd1 vccd1 vccd1 _5657_/X sky130_fd_sc_hd__buf_1
X_4608_ _7257_/Q _3899_/A _4616_/S vssd1 vssd1 vccd1 vccd1 _4609_/A sky130_fd_sc_hd__mux2_1
X_5588_ _5588_/A _6234_/C _6233_/B vssd1 vssd1 vccd1 vccd1 _5588_/X sky130_fd_sc_hd__or3_1
X_4539_ _4539_/A vssd1 vssd1 vccd1 vccd1 _7287_/D sky130_fd_sc_hd__clkbuf_1
X_7327_ _7525_/CLK _7327_/D vssd1 vssd1 vccd1 vccd1 _7327_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7258_ _7258_/CLK _7258_/D vssd1 vssd1 vccd1 vccd1 _7258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7189_ _7190_/CLK _7189_/D vssd1 vssd1 vccd1 vccd1 _7189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3083_ clkbuf_0__3083_/X vssd1 vssd1 vccd1 vccd1 _6320_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3910_ _3910_/A vssd1 vssd1 vccd1 vccd1 _7555_/D sky130_fd_sc_hd__clkbuf_1
X_4890_ _4831_/X _7076_/Q _4892_/S vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__mux2_1
X_3841_ _3841_/A vssd1 vssd1 vccd1 vccd1 _7582_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__3419_ clkbuf_0__3419_/X vssd1 vssd1 vccd1 vccd1 _6948__37/A sky130_fd_sc_hd__clkbuf_16
X_3772_ _3664_/X _7607_/Q _3774_/S vssd1 vssd1 vccd1 vccd1 _3773_/A sky130_fd_sc_hd__mux2_1
X_6560_ _6576_/D _6560_/B _6583_/C vssd1 vssd1 vccd1 vccd1 _6560_/X sky130_fd_sc_hd__and3b_1
XFILLER_9_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5511_ _6993_/A vssd1 vssd1 vccd1 vccd1 _7034_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6491_ _6482_/X _6483_/Y _6485_/X _6486_/Y _6490_/X vssd1 vssd1 vccd1 vccd1 _6491_/X
+ sky130_fd_sc_hd__a221o_1
X_5442_ _7724_/Q vssd1 vssd1 vccd1 vccd1 _6481_/A sky130_fd_sc_hd__buf_4
X_5373_ _5373_/A _5373_/B vssd1 vssd1 vccd1 vccd1 _5374_/A sky130_fd_sc_hd__or2_1
X_7112_ _7112_/CLK _7112_/D vssd1 vssd1 vccd1 vccd1 _7112_/Q sky130_fd_sc_hd__dfxtp_1
X_4324_ _4324_/A vssd1 vssd1 vccd1 vccd1 _7367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7043_ _7043_/CLK _7043_/D vssd1 vssd1 vccd1 vccd1 _7043_/Q sky130_fd_sc_hd__dfxtp_2
X_4255_ _7669_/Q vssd1 vssd1 vccd1 vccd1 _4255_/X sky130_fd_sc_hd__clkbuf_2
X_4186_ _4186_/A vssd1 vssd1 vccd1 vccd1 _7419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__2955_ _6031_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2955_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6827_ _6868_/A _6827_/B _6827_/C vssd1 vssd1 vccd1 vccd1 _6828_/A sky130_fd_sc_hd__and3_1
XFILLER_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6689_ _6713_/A vssd1 vssd1 vccd1 vccd1 _6689_/X sky130_fd_sc_hd__buf_1
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__2721_ clkbuf_0__2721_/X vssd1 vssd1 vccd1 vccd1 _5730__279/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3280_ clkbuf_0__3280_/X vssd1 vssd1 vccd1 vccd1 _6694__134/A sky130_fd_sc_hd__clkbuf_16
XFILLER_10_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4040_ _4936_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _4056_/S sky130_fd_sc_hd__nand2_2
Xclkbuf_4_12_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7525_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5991_ _6599_/A vssd1 vssd1 vccd1 vccd1 _5991_/X sky130_fd_sc_hd__clkbuf_2
X_4942_ _3804_/X _7041_/Q _4946_/S vssd1 vssd1 vccd1 vccd1 _4943_/A sky130_fd_sc_hd__mux2_1
X_7730_ _7731_/CLK _7730_/D vssd1 vssd1 vccd1 vccd1 _7730_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7661_ _7727_/CLK _7661_/D vssd1 vssd1 vccd1 vccd1 _7661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4873_ _4873_/A vssd1 vssd1 vccd1 vccd1 _7110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6612_ _7514_/Q _6609_/X _6611_/X _6569_/A vssd1 vssd1 vccd1 vccd1 _7514_/D sky130_fd_sc_hd__o211a_1
X_7592_ _7592_/CLK _7592_/D vssd1 vssd1 vccd1 vccd1 _7592_/Q sky130_fd_sc_hd__dfxtp_1
X_3824_ _4239_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _3840_/S sky130_fd_sc_hd__or2_4
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3755_ _3755_/A vssd1 vssd1 vccd1 vccd1 _7614_/D sky130_fd_sc_hd__clkbuf_1
X_6543_ _7501_/Q _6543_/B vssd1 vssd1 vccd1 vccd1 _6544_/C sky130_fd_sc_hd__or2_1
X_3686_ _3542_/X _7676_/Q _3688_/S vssd1 vssd1 vccd1 vccd1 _3687_/A sky130_fd_sc_hd__mux2_1
X_6474_ _7503_/Q _6474_/B _6474_/C vssd1 vssd1 vccd1 vccd1 _6474_/X sky130_fd_sc_hd__and3_1
X_5425_ _7533_/Q _7113_/Q _7565_/Q _7129_/Q _5252_/A _5138_/X vssd1 vssd1 vccd1 vccd1
+ _5425_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5356_ _5356_/A _5356_/B vssd1 vssd1 vccd1 vccd1 _5356_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_5 _3819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5287_ _5291_/A _5284_/Y _5286_/Y _5396_/A vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__o211a_1
X_4307_ _4307_/A vssd1 vssd1 vccd1 vccd1 _7374_/D sky130_fd_sc_hd__clkbuf_1
X_4238_ _7674_/Q vssd1 vssd1 vccd1 vccd1 _4238_/X sky130_fd_sc_hd__buf_4
Xclkbuf_0__3085_ _6302_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3085_/X sky130_fd_sc_hd__clkbuf_16
X_7026_ _7026_/A vssd1 vssd1 vccd1 vccd1 _7729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4169_ _4112_/X _7426_/Q _4173_/S vssd1 vssd1 vccd1 vccd1 _4170_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6435__66 _6437__68/A vssd1 vssd1 vccd1 vccd1 _7488_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6363__489 _6363__489/A vssd1 vssd1 vccd1 vccd1 _7431_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3540_ _3540_/A vssd1 vssd1 vccd1 vccd1 _7709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3471_ _7317_/Q vssd1 vssd1 vccd1 vccd1 _3900_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5210_ _5210_/A vssd1 vssd1 vccd1 vccd1 _5363_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5141_ _7542_/Q _7432_/Q _7400_/Q _7384_/Q _5138_/X _5293_/A vssd1 vssd1 vccd1 vccd1
+ _5141_/X sky130_fd_sc_hd__mux4_1
X_5072_ _5072_/A vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4023_ _3899_/X _7487_/Q _4031_/S vssd1 vssd1 vccd1 vccd1 _4024_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5974_ _7588_/Q _7580_/Q _7572_/Q _7486_/Q _5912_/X _5908_/X vssd1 vssd1 vccd1 vccd1
+ _5974_/X sky130_fd_sc_hd__mux4_2
XFILLER_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7713_ _7713_/CLK _7713_/D vssd1 vssd1 vccd1 vccd1 _7713_/Q sky130_fd_sc_hd__dfxtp_1
X_4925_ _4925_/A vssd1 vssd1 vccd1 vccd1 _7050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2723_ _5737_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2723_/X sky130_fd_sc_hd__clkbuf_16
X_4856_ _4834_/X _7117_/Q _4856_/S vssd1 vssd1 vccd1 vccd1 _4857_/A sky130_fd_sc_hd__mux2_1
X_7644_ _7655_/CLK _7644_/D vssd1 vssd1 vccd1 vccd1 _7644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7575_ _7575_/CLK _7575_/D vssd1 vssd1 vccd1 vccd1 _7575_/Q sky130_fd_sc_hd__dfxtp_1
X_3807_ _7671_/Q vssd1 vssd1 vccd1 vccd1 _3807_/X sky130_fd_sc_hd__buf_4
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6526_ _6524_/Y _6593_/C _6567_/A _6609_/A vssd1 vssd1 vccd1 vccd1 _6526_/X sky130_fd_sc_hd__a22o_1
X_4787_ _4787_/A vssd1 vssd1 vccd1 vccd1 _7145_/D sky130_fd_sc_hd__clkbuf_1
X_3738_ _3908_/A vssd1 vssd1 vccd1 vccd1 _3738_/X sky130_fd_sc_hd__buf_2
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3669_ _3668_/X _7683_/Q _3669_/S vssd1 vssd1 vccd1 vccd1 _3670_/A sky130_fd_sc_hd__mux2_1
X_6457_ _7511_/Q _6457_/B vssd1 vssd1 vccd1 vccd1 _6460_/A sky130_fd_sc_hd__xnor2_1
X_6388_ _6388_/A vssd1 vssd1 vccd1 vccd1 _6388_/X sky130_fd_sc_hd__buf_1
X_5408_ _7726_/Q vssd1 vssd1 vccd1 vccd1 _6133_/A sky130_fd_sc_hd__buf_4
XFILLER_87_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5339_ _5584_/B _5339_/B vssd1 vssd1 vccd1 vccd1 _5339_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7009_ _7009_/A vssd1 vssd1 vccd1 vccd1 _7724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4581_/X _7179_/Q _4712_/S vssd1 vssd1 vccd1 vccd1 _4711_/A sky130_fd_sc_hd__mux2_1
X_4641_ _4641_/A vssd1 vssd1 vccd1 vccd1 _7242_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4572_ _4572_/A vssd1 vssd1 vccd1 vccd1 _4572_/X sky130_fd_sc_hd__clkbuf_4
X_7360_ _7360_/CLK _7360_/D vssd1 vssd1 vccd1 vccd1 _7360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3523_ _3522_/X _7713_/Q _3535_/S vssd1 vssd1 vccd1 vccd1 _3524_/A sky130_fd_sc_hd__mux2_1
X_7291_ _7291_/CLK _7291_/D vssd1 vssd1 vccd1 vccd1 _7291_/Q sky130_fd_sc_hd__dfxtp_1
X_6242_ _6254_/A vssd1 vssd1 vccd1 vccd1 _6242_/X sky130_fd_sc_hd__buf_1
X_5659__221 _5661__223/A vssd1 vssd1 vccd1 vccd1 _7115_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5124_ _7095_/Q _7098_/Q _7102_/Q vssd1 vssd1 vccd1 vccd1 _5125_/D sky130_fd_sc_hd__or3_1
X_5055_ _5055_/A _5057_/B vssd1 vssd1 vccd1 vccd1 _5056_/A sky130_fd_sc_hd__and2_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4006_ _4006_/A vssd1 vssd1 vccd1 vccd1 _7495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5957_ _7247_/Q _7231_/Q _7477_/Q _7469_/Q _5925_/A _5861_/X vssd1 vssd1 vccd1 vccd1
+ _5957_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4908_ _4831_/X _7057_/Q _4910_/S vssd1 vssd1 vccd1 vccd1 _4909_/A sky130_fd_sc_hd__mux2_1
X_7627_ _7627_/CLK _7627_/D vssd1 vssd1 vccd1 vccd1 _7627_/Q sky130_fd_sc_hd__dfxtp_1
X_5888_ _5888_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5888_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4839_ _4839_/A vssd1 vssd1 vccd1 vccd1 _7124_/D sky130_fd_sc_hd__clkbuf_1
X_7558_ _7558_/CLK _7558_/D vssd1 vssd1 vccd1 vccd1 _7558_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_0__2637_ _5524_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2637_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7489_ _7489_/CLK _7489_/D vssd1 vssd1 vccd1 vccd1 _7489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6509_ _6509_/A _6509_/B _6509_/C _6508_/Y vssd1 vssd1 vccd1 vccd1 _6509_/X sky130_fd_sc_hd__or4b_1
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3100_ clkbuf_0__3100_/X vssd1 vssd1 vccd1 vccd1 _6385__507/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5504__184 _5504__184/A vssd1 vssd1 vccd1 vccd1 _7040_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6860_ _6860_/A vssd1 vssd1 vccd1 vccd1 _7651_/D sky130_fd_sc_hd__clkbuf_1
X_6791_ _6791_/A _6791_/B _6791_/C _6161_/B vssd1 vssd1 vccd1 vccd1 _6791_/X sky130_fd_sc_hd__or4b_1
X_5811_ _7497_/Q _7496_/Q vssd1 vssd1 vccd1 vccd1 _6607_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4624_ _4678_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _4640_/S sky130_fd_sc_hd__nand2_2
X_7412_ _7412_/CLK _7412_/D vssd1 vssd1 vccd1 vccd1 _7412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4555_ _4555_/A vssd1 vssd1 vccd1 vccd1 _7279_/D sky130_fd_sc_hd__clkbuf_1
X_7343_ _7343_/CLK _7343_/D vssd1 vssd1 vccd1 vccd1 _7343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3506_ _5645_/B _5123_/D _3506_/C _3506_/D vssd1 vssd1 vccd1 vccd1 _5586_/C sky130_fd_sc_hd__or4_4
X_4486_ _4477_/B _4486_/B _4486_/C vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__and3b_1
X_7274_ _7359_/CLK _7274_/D vssd1 vssd1 vccd1 vccd1 _7274_/Q sky130_fd_sc_hd__dfxtp_1
X_6225_ _7663_/Q _6231_/B vssd1 vssd1 vccd1 vccd1 _6226_/A sky130_fd_sc_hd__and2_1
XFILLER_112_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6474_/B _6791_/B vssd1 vssd1 vccd1 vccd1 _6774_/A sky130_fd_sc_hd__xnor2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5107_/A vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6249__400 _6253__404/A vssd1 vssd1 vccd1 vccd1 _7340_/CLK sky130_fd_sc_hd__inv_2
X_5038_ _5038_/A _5046_/B vssd1 vssd1 vccd1 vccd1 _5039_/A sky130_fd_sc_hd__and2_1
XFILLER_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6989_ _6989_/A vssd1 vssd1 vccd1 vccd1 _7718_/D sky130_fd_sc_hd__clkbuf_1
X_6952__40 _6956__44/A vssd1 vssd1 vccd1 vccd1 _7696_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2952_ clkbuf_0__2952_/X vssd1 vssd1 vccd1 vccd1 _6023__309/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput98 _5078_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[14] sky130_fd_sc_hd__buf_2
XFILLER_95_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_226 vssd1 vssd1 vccd1 vccd1 CaravelHost_226/HI versionID[0] sky130_fd_sc_hd__conb_1
XCaravelHost_215 vssd1 vssd1 vccd1 vccd1 CaravelHost_215/HI manufacturerID[7] sky130_fd_sc_hd__conb_1
XCaravelHost_204 vssd1 vssd1 vccd1 vccd1 CaravelHost_204/HI core1Index[4] sky130_fd_sc_hd__conb_1
XCaravelHost_237 vssd1 vssd1 vccd1 vccd1 partID[11] CaravelHost_237/LO sky130_fd_sc_hd__conb_1
X_4340_ _7322_/Q vssd1 vssd1 vccd1 vccd1 _4340_/X sky130_fd_sc_hd__clkbuf_4
X_4271_ _7389_/Q _3588_/X _4275_/S vssd1 vssd1 vccd1 vccd1 _4272_/A sky130_fd_sc_hd__mux2_1
X_6010_ _5902_/A _5999_/X _6009_/Y vssd1 vssd1 vccd1 vccd1 _6010_/X sky130_fd_sc_hd__a21o_1
X_6708__145 _6710__147/A vssd1 vssd1 vccd1 vccd1 _7589_/CLK sky130_fd_sc_hd__inv_2
X_6053__333 _6054__334/A vssd1 vssd1 vccd1 vccd1 _7259_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6912_ _6912_/A vssd1 vssd1 vccd1 vccd1 _7668_/D sky130_fd_sc_hd__clkbuf_1
X_6843_ _7648_/Q _6847_/C _6843_/C vssd1 vssd1 vccd1 vccd1 _6849_/B sky130_fd_sc_hd__and3_1
X_6631__83 _6632__84/A vssd1 vssd1 vccd1 vccd1 _7527_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3986_ _3633_/X _7524_/Q _3994_/S vssd1 vssd1 vccd1 vccd1 _3987_/A sky130_fd_sc_hd__mux2_1
X_6774_ _6774_/A _6774_/B _6774_/C _6774_/D vssd1 vssd1 vccd1 vccd1 _6779_/B sky130_fd_sc_hd__or4_1
XFILLER_22_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5725_ _5725_/A vssd1 vssd1 vccd1 vccd1 _5725_/X sky130_fd_sc_hd__buf_1
XFILLER_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6244__396 _6247__399/A vssd1 vssd1 vccd1 vccd1 _7336_/CLK sky130_fd_sc_hd__inv_2
X_4607_ _4622_/S vssd1 vssd1 vccd1 vccd1 _4616_/S sky130_fd_sc_hd__clkbuf_2
X_5587_ _5587_/A _5587_/B _5587_/C _5587_/D vssd1 vssd1 vccd1 vccd1 _6233_/B sky130_fd_sc_hd__or4_2
XFILLER_117_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4538_ _4232_/X _7287_/Q _4540_/S vssd1 vssd1 vccd1 vccd1 _4539_/A sky130_fd_sc_hd__mux2_1
X_7326_ _7525_/CLK _7326_/D vssd1 vssd1 vccd1 vccd1 _7326_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_116_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7257_ _7257_/CLK _7257_/D vssd1 vssd1 vccd1 vccd1 _7257_/Q sky130_fd_sc_hd__dfxtp_1
X_4469_ _5923_/A _4477_/A _4477_/B vssd1 vssd1 vccd1 vccd1 _4473_/B sky130_fd_sc_hd__and3_1
X_5704__258 _5705__259/A vssd1 vssd1 vccd1 vccd1 _7152_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6208_ _6214_/A vssd1 vssd1 vccd1 vccd1 _6208_/X sky130_fd_sc_hd__buf_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7188_ _7190_/CLK _7188_/D vssd1 vssd1 vccd1 vccd1 _7188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6139_ _6450_/B _6139_/B _6790_/A vssd1 vssd1 vccd1 vccd1 _6775_/B sky130_fd_sc_hd__and3_1
XFILLER_18_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3082_ clkbuf_0__3082_/X vssd1 vssd1 vccd1 vccd1 _6294__434/A sky130_fd_sc_hd__clkbuf_16
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3840_ _3753_/X _7582_/Q _3840_/S vssd1 vssd1 vccd1 vccd1 _3841_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__3418_ clkbuf_0__3418_/X vssd1 vssd1 vccd1 vccd1 _6944__34/A sky130_fd_sc_hd__clkbuf_16
X_3771_ _3771_/A vssd1 vssd1 vccd1 vccd1 _7608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5510_ _5535_/B vssd1 vssd1 vccd1 vccd1 _6993_/A sky130_fd_sc_hd__buf_2
XFILLER_118_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6490_ _6487_/X _6488_/X _6490_/S vssd1 vssd1 vccd1 vccd1 _6490_/X sky130_fd_sc_hd__mux2_1
X_5441_ _5469_/A _7275_/Q _6234_/B _5441_/D vssd1 vssd1 vccd1 vccd1 _5449_/A sky130_fd_sc_hd__and4_2
X_5372_ _6450_/A _5236_/A _5370_/Y _5371_/X _5112_/A vssd1 vssd1 vccd1 vccd1 _5373_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7111_ _7111_/CLK _7111_/D vssd1 vssd1 vccd1 vccd1 _7111_/Q sky130_fd_sc_hd__dfxtp_1
X_4323_ _7367_/Q _4320_/X _4335_/S vssd1 vssd1 vccd1 vccd1 _4324_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7042_ _7042_/CLK _7042_/D vssd1 vssd1 vccd1 vccd1 _7042_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4254_ _4254_/A vssd1 vssd1 vccd1 vccd1 _7395_/D sky130_fd_sc_hd__clkbuf_1
X_6680__123 _6680__123/A vssd1 vssd1 vccd1 vccd1 _7567_/CLK sky130_fd_sc_hd__inv_2
X_4185_ _4109_/X _7419_/Q _4185_/S vssd1 vssd1 vccd1 vccd1 _4186_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__2954_ _6025_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2954_/X sky130_fd_sc_hd__clkbuf_16
X_6826_ _6833_/C _6829_/C vssd1 vssd1 vccd1 vccd1 _6827_/C sky130_fd_sc_hd__or2_1
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6757_ _6763_/A vssd1 vssd1 vccd1 vccd1 _6757_/X sky130_fd_sc_hd__buf_1
XFILLER_50_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5710__262 _5712__264/A vssd1 vssd1 vccd1 vccd1 _7156_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3969_ _3644_/X _7532_/Q _3975_/S vssd1 vssd1 vccd1 vccd1 _3970_/A sky130_fd_sc_hd__mux2_1
X_6688_ _6688_/A vssd1 vssd1 vccd1 vccd1 _6688_/X sky130_fd_sc_hd__buf_1
X_5639_ _5639_/A vssd1 vssd1 vccd1 vccd1 _7101_/D sky130_fd_sc_hd__clkbuf_1
X_7309_ _7309_/CLK _7309_/D vssd1 vssd1 vccd1 vccd1 _7309_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__2720_ clkbuf_0__2720_/X vssd1 vssd1 vccd1 vccd1 _5724__274/A sky130_fd_sc_hd__clkbuf_16
XFILLER_86_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5653__216 _5656__219/A vssd1 vssd1 vccd1 vccd1 _7110_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5990_ _5882_/X _5979_/X _5989_/Y vssd1 vssd1 vccd1 vccd1 _5990_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4941_ _4941_/A vssd1 vssd1 vccd1 vccd1 _7042_/D sky130_fd_sc_hd__clkbuf_1
X_7660_ _7727_/CLK _7660_/D vssd1 vssd1 vccd1 vccd1 _7660_/Q sky130_fd_sc_hd__dfxtp_1
X_4872_ _4831_/X _7110_/Q _4874_/S vssd1 vssd1 vccd1 vccd1 _4873_/A sky130_fd_sc_hd__mux2_1
X_3823_ _4095_/B _3900_/C _4095_/A vssd1 vssd1 vccd1 vccd1 _4021_/B sky130_fd_sc_hd__or3b_4
X_6611_ _7516_/Q _7515_/Q _6609_/A _6593_/C _6610_/Y vssd1 vssd1 vccd1 vccd1 _6611_/X
+ sky130_fd_sc_hd__a311o_1
X_7591_ _7591_/CLK _7591_/D vssd1 vssd1 vccd1 vccd1 _7591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3754_ _3753_/X _7614_/Q _3754_/S vssd1 vssd1 vccd1 vccd1 _3755_/A sky130_fd_sc_hd__mux2_1
X_6542_ _6558_/D vssd1 vssd1 vccd1 vccd1 _6553_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3685_ _3685_/A vssd1 vssd1 vccd1 vccd1 _7677_/D sky130_fd_sc_hd__clkbuf_1
X_6473_ _6474_/B _6474_/C _6558_/B vssd1 vssd1 vccd1 vccd1 _6473_/Y sky130_fd_sc_hd__a21oi_1
X_5424_ _5365_/A _5423_/X _5213_/A vssd1 vssd1 vccd1 vccd1 _5424_/X sky130_fd_sc_hd__a21o_1
X_5355_ _7531_/Q _7111_/Q _7563_/Q _7127_/Q _5132_/X _5135_/X vssd1 vssd1 vccd1 vccd1
+ _5356_/B sky130_fd_sc_hd__mux4_1
XINSDIODE2_6 _3911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4306_ _4217_/X _7374_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4307_/A sky130_fd_sc_hd__mux2_1
X_5286_ _5360_/A _5286_/B vssd1 vssd1 vccd1 vccd1 _5286_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3084_ _6296_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3084_/X sky130_fd_sc_hd__clkbuf_16
X_4237_ _4237_/A vssd1 vssd1 vccd1 vccd1 _7400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7025_ _7031_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _7026_/A sky130_fd_sc_hd__and2b_1
XFILLER_114_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4168_ _4168_/A vssd1 vssd1 vccd1 vccd1 _7427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4099_ _4099_/A vssd1 vssd1 vccd1 vccd1 _7455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6066__343 _6067__344/A vssd1 vssd1 vccd1 vccd1 _7269_/CLK sky130_fd_sc_hd__inv_2
X_6809_ _6809_/A vssd1 vssd1 vccd1 vccd1 _6859_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6687__129 _6687__129/A vssd1 vssd1 vccd1 vccd1 _7573_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5717__268 _5718__269/A vssd1 vssd1 vccd1 vccd1 _7162_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3470_ _7319_/Q vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5140_ _5148_/A vssd1 vssd1 vccd1 vccd1 _5293_/A sky130_fd_sc_hd__buf_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5071_ _5071_/A _5079_/B vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__and2_1
XFILLER_96_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4022_ _4037_/S vssd1 vssd1 vccd1 vccd1 _4031_/S sky130_fd_sc_hd__buf_2
XFILLER_77_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5973_ _7540_/Q _7681_/Q _7697_/Q _7283_/Q _5907_/X _5905_/X vssd1 vssd1 vccd1 vccd1
+ _5973_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7712_ _7712_/CLK _7712_/D vssd1 vssd1 vccd1 vccd1 _7712_/Q sky130_fd_sc_hd__dfxtp_1
X_4924_ _7050_/Q _4569_/A _4928_/S vssd1 vssd1 vccd1 vccd1 _4925_/A sky130_fd_sc_hd__mux2_1
X_6440__70 _6441__71/A vssd1 vssd1 vccd1 vccd1 _7492_/CLK sky130_fd_sc_hd__inv_2
X_4855_ _4855_/A vssd1 vssd1 vccd1 vccd1 _7118_/D sky130_fd_sc_hd__clkbuf_1
X_7643_ _7655_/CLK _7643_/D vssd1 vssd1 vccd1 vccd1 _7643_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2722_ _5731_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2722_/X sky130_fd_sc_hd__clkbuf_16
X_7574_ _7574_/CLK _7574_/D vssd1 vssd1 vccd1 vccd1 _7574_/Q sky130_fd_sc_hd__dfxtp_1
X_3806_ _3806_/A vssd1 vssd1 vccd1 vccd1 _7595_/D sky130_fd_sc_hd__clkbuf_1
X_4786_ _7145_/Q _4560_/A _4794_/S vssd1 vssd1 vccd1 vccd1 _4787_/A sky130_fd_sc_hd__mux2_1
X_3737_ _3737_/A vssd1 vssd1 vccd1 vccd1 _7620_/D sky130_fd_sc_hd__clkbuf_1
X_6525_ _6525_/A vssd1 vssd1 vccd1 vccd1 _6593_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3668_ _4584_/A vssd1 vssd1 vccd1 vccd1 _3668_/X sky130_fd_sc_hd__buf_2
X_6456_ _7718_/Q _6107_/A _6112_/A vssd1 vssd1 vccd1 vccd1 _6457_/B sky130_fd_sc_hd__a21oi_1
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3599_ _3599_/A vssd1 vssd1 vccd1 vccd1 _7701_/D sky130_fd_sc_hd__clkbuf_1
X_5407_ _4384_/A _5396_/X _5400_/X _5406_/X _5433_/A vssd1 vssd1 vccd1 vccd1 _5407_/X
+ sky130_fd_sc_hd__a311o_1
X_5338_ _5161_/X _5322_/X _5337_/X _5308_/A vssd1 vssd1 vccd1 vccd1 _5338_/X sky130_fd_sc_hd__a211o_1
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7008_ _7003_/X _7008_/B vssd1 vssd1 vccd1 vccd1 _7009_/A sky130_fd_sc_hd__and2b_1
X_5269_ _5365_/A _5268_/X vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__or2b_1
XFILLER_56_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6959__46 _6962__49/A vssd1 vssd1 vccd1 vccd1 _7702_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6693__133 _6694__134/A vssd1 vssd1 vccd1 vccd1 _7577_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4640_ _4261_/X _7242_/Q _4640_/S vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4571_ _4571_/A vssd1 vssd1 vccd1 vccd1 _7271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3522_ _3905_/A vssd1 vssd1 vccd1 vccd1 _3522_/X sky130_fd_sc_hd__buf_2
X_7290_ _7290_/CLK _7290_/D vssd1 vssd1 vccd1 vccd1 _7290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6017__304 _6017__304/A vssd1 vssd1 vccd1 vccd1 _7230_/CLK sky130_fd_sc_hd__inv_2
X_5123_ _7099_/Q _7100_/Q _7101_/Q _5123_/D vssd1 vssd1 vccd1 vccd1 _5126_/C sky130_fd_sc_hd__or4_1
X_6638__89 _6638__89/A vssd1 vssd1 vccd1 vccd1 _7533_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5054_/A vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4005_ _7495_/Q _3549_/X _4013_/S vssd1 vssd1 vccd1 vccd1 _4006_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _5954_/X _5955_/X _5995_/S vssd1 vssd1 vccd1 vccd1 _5956_/X sky130_fd_sc_hd__mux2_2
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5887_ _7394_/Q _7236_/Q _7552_/Q _7458_/Q _5857_/X _4484_/X vssd1 vssd1 vccd1 vccd1
+ _5888_/B sky130_fd_sc_hd__mux4_1
X_4907_ _4907_/A vssd1 vssd1 vccd1 vccd1 _7058_/D sky130_fd_sc_hd__clkbuf_1
X_7626_ _7626_/CLK _7626_/D vssd1 vssd1 vccd1 vccd1 _7626_/Q sky130_fd_sc_hd__dfxtp_1
X_4838_ _4837_/X _7124_/Q _4844_/S vssd1 vssd1 vccd1 vccd1 _4839_/A sky130_fd_sc_hd__mux2_1
X_7557_ _7557_/CLK _7557_/D vssd1 vssd1 vccd1 vccd1 _7557_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2636_ _5518_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2636_/X sky130_fd_sc_hd__clkbuf_16
X_4769_ _4769_/A vssd1 vssd1 vccd1 vccd1 _7153_/D sky130_fd_sc_hd__clkbuf_1
X_7488_ _7488_/CLK _7488_/D vssd1 vssd1 vccd1 vccd1 _7488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6508_ _6485_/X _6486_/Y _6454_/D _6490_/X _6507_/X vssd1 vssd1 vccd1 vccd1 _6508_/Y
+ sky130_fd_sc_hd__a2111oi_1
X_6439_ _6619_/A vssd1 vssd1 vccd1 vccd1 _6439_/X sky130_fd_sc_hd__buf_1
XFILLER_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6790_ _6790_/A vssd1 vssd1 vccd1 vccd1 _6791_/A sky130_fd_sc_hd__clkinv_2
XFILLER_35_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7411_ _7411_/CLK _7411_/D vssd1 vssd1 vccd1 vccd1 _7411_/Q sky130_fd_sc_hd__dfxtp_1
X_4623_ _4623_/A vssd1 vssd1 vccd1 vccd1 _7250_/D sky130_fd_sc_hd__clkbuf_1
X_4554_ _7279_/Q _3917_/A _4558_/S vssd1 vssd1 vccd1 vccd1 _4555_/A sky130_fd_sc_hd__mux2_1
X_7342_ _7342_/CLK _7342_/D vssd1 vssd1 vccd1 vccd1 _7342_/Q sky130_fd_sc_hd__dfxtp_1
X_7273_ _7273_/CLK _7273_/D vssd1 vssd1 vccd1 vccd1 _7273_/Q sky130_fd_sc_hd__dfxtp_1
X_3505_ _7095_/Q _7096_/Q _7097_/Q _7098_/Q vssd1 vssd1 vccd1 vccd1 _3506_/D sky130_fd_sc_hd__or4_1
X_4485_ _7330_/Q _6236_/C _4484_/X vssd1 vssd1 vccd1 vccd1 _4486_/B sky130_fd_sc_hd__a21o_1
X_6224_ _6224_/A vssd1 vssd1 vccd1 vccd1 _7324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6476_/A _7646_/Q vssd1 vssd1 vccd1 vccd1 _6791_/B sky130_fd_sc_hd__xor2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _7205_/Q _5106_/B vssd1 vssd1 vccd1 vccd1 _5107_/A sky130_fd_sc_hd__and2_1
X_6086_ _6086_/A vssd1 vssd1 vccd1 vccd1 _6086_/X sky130_fd_sc_hd__buf_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5037_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5046_/B sky130_fd_sc_hd__buf_4
XFILLER_85_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6988_ _6981_/X _6988_/B vssd1 vssd1 vccd1 vccd1 _6989_/A sky130_fd_sc_hd__and2b_1
XFILLER_15_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5939_ _7246_/Q _7230_/Q _7476_/Q _7468_/Q _5860_/X _5861_/X vssd1 vssd1 vccd1 vccd1
+ _5939_/X sky130_fd_sc_hd__mux4_1
X_7609_ _7609_/CLK _7609_/D vssd1 vssd1 vccd1 vccd1 _7609_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2951_ clkbuf_0__2951_/X vssd1 vssd1 vccd1 vccd1 _6017__304/A sky130_fd_sc_hd__clkbuf_16
Xoutput99 _5080_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[15] sky130_fd_sc_hd__buf_2
XFILLER_103_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XCaravelHost_227 vssd1 vssd1 vccd1 vccd1 CaravelHost_227/HI versionID[1] sky130_fd_sc_hd__conb_1
XCaravelHost_216 vssd1 vssd1 vccd1 vccd1 CaravelHost_216/HI manufacturerID[8] sky130_fd_sc_hd__conb_1
XCaravelHost_205 vssd1 vssd1 vccd1 vccd1 CaravelHost_205/HI core1Index[5] sky130_fd_sc_hd__conb_1
XCaravelHost_238 vssd1 vssd1 vccd1 vccd1 partID[14] CaravelHost_238/LO sky130_fd_sc_hd__conb_1
XFILLER_99_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4270_ _4270_/A vssd1 vssd1 vccd1 vccd1 _7390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6911_ _6911_/A _6921_/B _6921_/C vssd1 vssd1 vccd1 vccd1 _6912_/A sky130_fd_sc_hd__and3_1
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6842_ _6842_/A vssd1 vssd1 vccd1 vccd1 _7647_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3985_ _4000_/S vssd1 vssd1 vccd1 vccd1 _3994_/S sky130_fd_sc_hd__buf_2
X_6773_ _6121_/Y _6122_/X _6126_/Y _6788_/A _6147_/Y vssd1 vssd1 vccd1 vccd1 _6774_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6060__338 _6060__338/A vssd1 vssd1 vccd1 vccd1 _7264_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4606_ _4606_/A _4606_/B _4936_/B vssd1 vssd1 vccd1 vccd1 _4622_/S sky130_fd_sc_hd__and3_2
X_5586_ _7089_/Q _7090_/Q _5586_/C vssd1 vssd1 vccd1 vccd1 _5587_/D sky130_fd_sc_hd__or3_1
X_7325_ _7525_/CLK _7325_/D vssd1 vssd1 vccd1 vccd1 _7325_/Q sky130_fd_sc_hd__dfxtp_4
X_4537_ _4537_/A vssd1 vssd1 vccd1 vccd1 _7288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7256_ _7256_/CLK _7256_/D vssd1 vssd1 vccd1 vccd1 _7256_/Q sky130_fd_sc_hd__dfxtp_1
X_4468_ _4468_/A _7330_/Q _4483_/A vssd1 vssd1 vccd1 vccd1 _4477_/B sky130_fd_sc_hd__and3_1
XFILLER_89_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6207_ _6207_/A vssd1 vssd1 vccd1 vccd1 _6207_/X sky130_fd_sc_hd__buf_1
X_7187_ _7190_/CLK _7187_/D vssd1 vssd1 vccd1 vccd1 _7187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6138_ _6483_/B _6139_/B _6790_/A vssd1 vssd1 vccd1 vccd1 _6775_/A sky130_fd_sc_hd__a21oi_1
X_4399_ _4399_/A vssd1 vssd1 vccd1 vccd1 _7347_/D sky130_fd_sc_hd__clkbuf_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3081_ clkbuf_0__3081_/X vssd1 vssd1 vccd1 vccd1 _6287__428/A sky130_fd_sc_hd__clkbuf_16
XFILLER_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6759__11 _6761__13/A vssd1 vssd1 vccd1 vccd1 _7630_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__3417_ clkbuf_0__3417_/X vssd1 vssd1 vccd1 vccd1 _6963_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3770_ _3660_/X _7608_/Q _3774_/S vssd1 vssd1 vccd1 vccd1 _3771_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__3279_ clkbuf_0__3279_/X vssd1 vssd1 vccd1 vccd1 _6713_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_13_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5440_ _5440_/A vssd1 vssd1 vccd1 vccd1 _6234_/B sky130_fd_sc_hd__clkbuf_2
X_6714__150 _6716__152/A vssd1 vssd1 vccd1 vccd1 _7594_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5371_ _7320_/Q _5339_/B _5469_/C vssd1 vssd1 vccd1 vccd1 _5371_/X sky130_fd_sc_hd__a21o_1
X_4322_ _4344_/S vssd1 vssd1 vccd1 vccd1 _4335_/S sky130_fd_sc_hd__buf_2
X_7110_ _7110_/CLK _7110_/D vssd1 vssd1 vccd1 vccd1 _7110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4253_ _4252_/X _7395_/Q _4253_/S vssd1 vssd1 vccd1 vccd1 _4254_/A sky130_fd_sc_hd__mux2_1
X_7041_ _7041_/CLK _7041_/D vssd1 vssd1 vccd1 vccd1 _7041_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4184_ _4184_/A vssd1 vssd1 vccd1 vccd1 _7420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2953_ _6024_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2953_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_63_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6825_ _6833_/C _6829_/C vssd1 vssd1 vccd1 vccd1 _6827_/B sky130_fd_sc_hd__nand2_1
X_3968_ _3968_/A vssd1 vssd1 vccd1 vccd1 _7533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5707_ _5731_/A vssd1 vssd1 vccd1 vccd1 _5707_/X sky130_fd_sc_hd__buf_1
X_3899_ _3899_/A vssd1 vssd1 vccd1 vccd1 _3899_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5638_ _7101_/Q _7200_/Q _6076_/S vssd1 vssd1 vccd1 vccd1 _5639_/A sky130_fd_sc_hd__mux2_1
X_5569_ _6561_/A vssd1 vssd1 vccd1 vccd1 _6609_/A sky130_fd_sc_hd__clkbuf_2
X_7308_ _7308_/CLK _7308_/D vssd1 vssd1 vccd1 vccd1 _7308_/Q sky130_fd_sc_hd__dfxtp_1
X_7239_ _7239_/CLK _7239_/D vssd1 vssd1 vccd1 vccd1 _7239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6269__415 _6276__419/A vssd1 vssd1 vccd1 vccd1 _7355_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4940_ _3801_/X _7042_/Q _4946_/S vssd1 vssd1 vccd1 vccd1 _4941_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4871_ _4871_/A vssd1 vssd1 vccd1 vccd1 _7111_/D sky130_fd_sc_hd__clkbuf_1
X_7590_ _7590_/CLK _7590_/D vssd1 vssd1 vccd1 vccd1 _7590_/Q sky130_fd_sc_hd__dfxtp_1
X_3822_ _3822_/A _6233_/A _3822_/C _3796_/C vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__or4b_4
XFILLER_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6610_ _7514_/Q _6610_/B vssd1 vssd1 vccd1 vccd1 _6610_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6541_ _7501_/Q _6541_/B _6541_/C _7498_/Q vssd1 vssd1 vccd1 vccd1 _6558_/D sky130_fd_sc_hd__and4_1
X_3753_ _3923_/A vssd1 vssd1 vccd1 vccd1 _3753_/X sky130_fd_sc_hd__buf_2
XFILLER_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3684_ _3538_/X _7677_/Q _3688_/S vssd1 vssd1 vccd1 vccd1 _3685_/A sky130_fd_sc_hd__mux2_1
X_6276__419 _6276__419/A vssd1 vssd1 vccd1 vccd1 _7361_/CLK sky130_fd_sc_hd__inv_2
X_6472_ _7503_/Q vssd1 vssd1 vccd1 vccd1 _6558_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5423_ _7690_/Q _7613_/Q _5429_/S vssd1 vssd1 vccd1 vccd1 _5423_/X sky130_fd_sc_hd__mux2_1
X_5354_ _5205_/X _5349_/X _5351_/Y _5353_/Y vssd1 vssd1 vccd1 vccd1 _5354_/X sky130_fd_sc_hd__o2bb2a_1
X_4305_ _4305_/A vssd1 vssd1 vccd1 vccd1 _7375_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_7 _3914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5285_ _7686_/Q _7609_/Q _5285_/S vssd1 vssd1 vccd1 vccd1 _5286_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3083_ _6295_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3083_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4236_ _4235_/X _7400_/Q _4236_/S vssd1 vssd1 vccd1 vccd1 _4237_/A sky130_fd_sc_hd__mux2_1
X_7024_ _6915_/A _5281_/X _7024_/S vssd1 vssd1 vccd1 vccd1 _7025_/B sky130_fd_sc_hd__mux2_1
X_4167_ _4109_/X _7427_/Q _4167_/S vssd1 vssd1 vccd1 vccd1 _4168_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4098_ _4094_/X _7455_/Q _4110_/S vssd1 vssd1 vccd1 vccd1 _4099_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6808_ _6808_/A vssd1 vssd1 vccd1 vccd1 _7640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3419_ _6945_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3419_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_105_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5572__204 _5572__204/A vssd1 vssd1 vccd1 vccd1 _7072_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5070_ _5092_/A vssd1 vssd1 vccd1 vccd1 _5079_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4021_ _4175_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _4037_/S sky130_fd_sc_hd__or2_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5972_ _7223_/Q _5814_/A _5971_/X _5880_/X vssd1 vssd1 vccd1 vccd1 _7223_/D sky130_fd_sc_hd__o211a_1
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7711_ _7711_/CLK _7711_/D vssd1 vssd1 vccd1 vccd1 _7711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4923_ _4923_/A vssd1 vssd1 vccd1 vccd1 _7051_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__2721_ _5725_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2721_/X sky130_fd_sc_hd__clkbuf_16
X_7642_ _7655_/CLK _7642_/D vssd1 vssd1 vccd1 vccd1 _7642_/Q sky130_fd_sc_hd__dfxtp_1
X_4854_ _4831_/X _7118_/Q _4856_/S vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7573_ _7573_/CLK _7573_/D vssd1 vssd1 vccd1 vccd1 _7573_/Q sky130_fd_sc_hd__dfxtp_1
X_3805_ _7595_/Q _3804_/X _3811_/S vssd1 vssd1 vccd1 vccd1 _3806_/A sky130_fd_sc_hd__mux2_1
X_4785_ _4800_/S vssd1 vssd1 vccd1 vccd1 _4794_/S sky130_fd_sc_hd__buf_2
X_3736_ _3735_/X _7620_/Q _3745_/S vssd1 vssd1 vccd1 vccd1 _3737_/A sky130_fd_sc_hd__mux2_1
X_6524_ _6532_/C vssd1 vssd1 vccd1 vccd1 _6524_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3667_ _7321_/Q vssd1 vssd1 vccd1 vccd1 _4584_/A sky130_fd_sc_hd__buf_2
X_6455_ _6504_/D _6455_/B vssd1 vssd1 vccd1 vccd1 _6572_/A sky130_fd_sc_hd__nor2_1
X_3598_ _7701_/Q _3597_/X _3604_/S vssd1 vssd1 vccd1 vccd1 _3599_/A sky130_fd_sc_hd__mux2_1
X_5406_ _5402_/X _5404_/X _5405_/X _5396_/A _5205_/A vssd1 vssd1 vccd1 vccd1 _5406_/X
+ sky130_fd_sc_hd__o221a_1
X_5337_ _5337_/A _5337_/B _5337_/C vssd1 vssd1 vccd1 vccd1 _5337_/X sky130_fd_sc_hd__and3_1
X_5268_ _7519_/Q _7140_/Q _5299_/A vssd1 vssd1 vccd1 vccd1 _5268_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4219_ _4219_/A vssd1 vssd1 vccd1 vccd1 _7406_/D sky130_fd_sc_hd__clkbuf_1
X_7007_ _4993_/A _6481_/A _7007_/S vssd1 vssd1 vccd1 vccd1 _7008_/B sky130_fd_sc_hd__mux2_1
X_6727__160 _6729__162/A vssd1 vssd1 vccd1 vccd1 _7604_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5199_ _5245_/A vssd1 vssd1 vccd1 vccd1 _5391_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5723__273 _5723__273/A vssd1 vssd1 vccd1 vccd1 _7167_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6346__475 _6347__476/A vssd1 vssd1 vccd1 vccd1 _7417_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4570_ _4569_/X _7271_/Q _4576_/S vssd1 vssd1 vccd1 vccd1 _4571_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3521_ _7673_/Q vssd1 vssd1 vccd1 vccd1 _3905_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6171_ _6171_/A vssd1 vssd1 vccd1 vccd1 _7285_/D sky130_fd_sc_hd__clkbuf_1
X_5122_ _5232_/A _5232_/B vssd1 vssd1 vccd1 vccd1 _5469_/C sky130_fd_sc_hd__nor2_2
XFILLER_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5053_ _5053_/A _5057_/B vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__and2_1
X_4004_ _4019_/S vssd1 vssd1 vccd1 vccd1 _4013_/S sky130_fd_sc_hd__clkbuf_2
X_5520__191 _5523__194/A vssd1 vssd1 vccd1 vccd1 _7048_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__2959_ clkbuf_0__2959_/X vssd1 vssd1 vccd1 vccd1 _6086_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_65_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5955_ _7587_/Q _7579_/Q _7571_/Q _7485_/Q _5912_/X _5908_/X vssd1 vssd1 vccd1 vccd1
+ _5955_/X sky130_fd_sc_hd__mux4_2
X_5886_ _5966_/A _5886_/B vssd1 vssd1 vccd1 vccd1 _5886_/Y sky130_fd_sc_hd__nor2_1
X_6964__50 _6967__53/A vssd1 vssd1 vccd1 vccd1 _7706_/CLK sky130_fd_sc_hd__inv_2
X_4906_ _4828_/X _7058_/Q _4910_/S vssd1 vssd1 vccd1 vccd1 _4907_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7625_ _7625_/CLK _7625_/D vssd1 vssd1 vccd1 vccd1 _7625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4837_ _7323_/Q vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5666__227 _5667__228/A vssd1 vssd1 vccd1 vccd1 _7121_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7556_ _7556_/CLK _7556_/D vssd1 vssd1 vccd1 vccd1 _7556_/Q sky130_fd_sc_hd__dfxtp_2
X_4768_ _7153_/Q _4320_/X _4774_/S vssd1 vssd1 vccd1 vccd1 _4769_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7487_ _7487_/CLK _7487_/D vssd1 vssd1 vccd1 vccd1 _7487_/Q sky130_fd_sc_hd__dfxtp_1
X_3719_ _3719_/A vssd1 vssd1 vccd1 vccd1 _7627_/D sky130_fd_sc_hd__clkbuf_1
X_4699_ _4699_/A vssd1 vssd1 vccd1 vccd1 _7185_/D sky130_fd_sc_hd__clkbuf_1
X_6507_ _7504_/Q _6507_/B _6507_/C vssd1 vssd1 vccd1 vccd1 _6507_/X sky130_fd_sc_hd__and3_1
XFILLER_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6643__93 _6644__94/A vssd1 vssd1 vccd1 vccd1 _7537_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7410_ _7410_/CLK _7410_/D vssd1 vssd1 vccd1 vccd1 _7410_/Q sky130_fd_sc_hd__dfxtp_1
X_4622_ _7250_/Q _3923_/A _4622_/S vssd1 vssd1 vccd1 vccd1 _4623_/A sky130_fd_sc_hd__mux2_1
X_4553_ _4553_/A vssd1 vssd1 vccd1 vccd1 _7280_/D sky130_fd_sc_hd__clkbuf_1
X_7341_ _7341_/CLK _7341_/D vssd1 vssd1 vccd1 vccd1 _7341_/Q sky130_fd_sc_hd__dfxtp_1
X_7272_ _7272_/CLK _7272_/D vssd1 vssd1 vccd1 vccd1 _7272_/Q sky130_fd_sc_hd__dfxtp_1
X_4484_ _5884_/A vssd1 vssd1 vccd1 vccd1 _4484_/X sky130_fd_sc_hd__buf_4
X_3504_ _7099_/Q _7100_/Q _7101_/Q _7102_/Q vssd1 vssd1 vccd1 vccd1 _3506_/C sky130_fd_sc_hd__or4_1
XFILLER_89_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6223_ _7662_/Q _6231_/B vssd1 vssd1 vccd1 vccd1 _6224_/A sky130_fd_sc_hd__and2_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3089_ clkbuf_0__3089_/X vssd1 vssd1 vccd1 vccd1 _6333_/A sky130_fd_sc_hd__clkbuf_16
X_6154_ _6483_/B _6483_/C vssd1 vssd1 vccd1 vccd1 _6474_/B sky130_fd_sc_hd__nand2_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5105_/A vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5036_/A vssd1 vssd1 vccd1 vccd1 _5036_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6987_ _5006_/A _7718_/Q _7000_/S vssd1 vssd1 vccd1 vccd1 _6988_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5938_ _7214_/Q _7040_/Q _7262_/Q _7254_/Q _5912_/X _5913_/X vssd1 vssd1 vccd1 vccd1
+ _5938_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5869_ _5869_/A vssd1 vssd1 vccd1 vccd1 _5998_/S sky130_fd_sc_hd__clkbuf_2
X_7608_ _7608_/CLK _7608_/D vssd1 vssd1 vccd1 vccd1 _7608_/Q sky130_fd_sc_hd__dfxtp_1
X_7539_ _7539_/CLK _7539_/D vssd1 vssd1 vccd1 vccd1 _7539_/Q sky130_fd_sc_hd__dfxtp_1
X_6256__406 _6256__406/A vssd1 vssd1 vccd1 vccd1 _7346_/CLK sky130_fd_sc_hd__inv_2
X_5527__197 _5529__199/A vssd1 vssd1 vccd1 vccd1 _7054_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XCaravelHost_217 vssd1 vssd1 vccd1 vccd1 CaravelHost_217/HI manufacturerID[9] sky130_fd_sc_hd__conb_1
XCaravelHost_206 vssd1 vssd1 vccd1 vccd1 CaravelHost_206/HI core1Index[6] sky130_fd_sc_hd__conb_1
XCaravelHost_228 vssd1 vssd1 vccd1 vccd1 CaravelHost_228/HI versionID[2] sky130_fd_sc_hd__conb_1
XCaravelHost_239 vssd1 vssd1 vccd1 vccd1 partID[15] CaravelHost_239/LO sky130_fd_sc_hd__conb_1
X_6196__375 _6199__378/A vssd1 vssd1 vccd1 vccd1 _7305_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_9_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7727_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_79_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6910_ _3511_/A _6910_/B vssd1 vssd1 vccd1 vccd1 _6921_/B sky130_fd_sc_hd__and2b_2
XFILLER_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6841_ _6868_/A _6841_/B _6841_/C vssd1 vssd1 vccd1 vccd1 _6842_/A sky130_fd_sc_hd__and3_1
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6402__520 _6403__521/A vssd1 vssd1 vccd1 vccd1 _7462_/CLK sky130_fd_sc_hd__inv_2
X_3984_ _4802_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _4000_/S sky130_fd_sc_hd__or2_2
X_6772_ _6134_/Y _6135_/X _6143_/Y _6131_/X vssd1 vssd1 vccd1 vccd1 _6774_/C sky130_fd_sc_hd__a211o_1
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4605_ _4605_/A vssd1 vssd1 vccd1 vccd1 _7258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6359__485 _6360__486/A vssd1 vssd1 vccd1 vccd1 _7427_/CLK sky130_fd_sc_hd__inv_2
X_5585_ _7082_/Q _5585_/B _5585_/C vssd1 vssd1 vccd1 vccd1 _5587_/A sky130_fd_sc_hd__or3_1
X_7324_ _7727_/CLK _7324_/D vssd1 vssd1 vccd1 vccd1 _7324_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4536_ _4229_/X _7288_/Q _4540_/S vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__mux2_1
X_7255_ _7255_/CLK _7255_/D vssd1 vssd1 vccd1 vccd1 _7255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4467_ _3484_/B _4467_/B _4467_/C vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__nand3b_1
XFILLER_98_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7186_ _7190_/CLK _7186_/D vssd1 vssd1 vccd1 vccd1 _7186_/Q sky130_fd_sc_hd__dfxtp_1
X_4398_ _4393_/B _4398_/B _6272_/C vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__and3b_1
X_6137_ _6137_/A _7648_/Q vssd1 vssd1 vccd1 vccd1 _6790_/A sky130_fd_sc_hd__xnor2_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6068_ _6086_/A vssd1 vssd1 vccd1 vccd1 _6068_/X sky130_fd_sc_hd__buf_1
X_5019_ _5019_/A vssd1 vssd1 vccd1 vccd1 _5019_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6303__440 _6304__441/A vssd1 vssd1 vccd1 vccd1 _7382_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3080_ clkbuf_0__3080_/X vssd1 vssd1 vccd1 vccd1 _6281__423/A sky130_fd_sc_hd__clkbuf_16
XFILLER_107_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5679__237 _5679__237/A vssd1 vssd1 vccd1 vccd1 _7131_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__3416_ clkbuf_0__3416_/X vssd1 vssd1 vccd1 vccd1 _6934__26/A sky130_fd_sc_hd__clkbuf_16
XFILLER_83_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__3278_ clkbuf_0__3278_/X vssd1 vssd1 vccd1 vccd1 _6687__129/A sky130_fd_sc_hd__clkbuf_16
XFILLER_80_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6204__382 _6204__382/A vssd1 vssd1 vccd1 vccd1 _7312_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5370_ _5337_/A _5354_/X _5369_/X _5308_/A vssd1 vssd1 vccd1 vccd1 _5370_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4321_ _4882_/A _4562_/A vssd1 vssd1 vccd1 vccd1 _4344_/S sky130_fd_sc_hd__nor2_2
X_7040_ _7040_/CLK _7040_/D vssd1 vssd1 vccd1 vccd1 _7040_/Q sky130_fd_sc_hd__dfxtp_1
X_4252_ _7670_/Q vssd1 vssd1 vccd1 vccd1 _4252_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4183_ _4106_/X _7420_/Q _4185_/S vssd1 vssd1 vccd1 vccd1 _4184_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6721__155 _6724__158/A vssd1 vssd1 vccd1 vccd1 _7599_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__2952_ _6018_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2952_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6824_ _7644_/Q vssd1 vssd1 vccd1 vccd1 _6833_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3967_ _3633_/X _7533_/Q _3975_/S vssd1 vssd1 vccd1 vccd1 _3968_/A sky130_fd_sc_hd__mux2_1
X_5706_ _5706_/A vssd1 vssd1 vccd1 vccd1 _5706_/X sky130_fd_sc_hd__buf_1
X_3898_ _3898_/A vssd1 vssd1 vccd1 vccd1 _7558_/D sky130_fd_sc_hd__clkbuf_1
X_5637_ _5637_/A vssd1 vssd1 vccd1 vccd1 _6076_/S sky130_fd_sc_hd__buf_4
XFILLER_88_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5568_ _5566_/X _5567_/X _7516_/Q vssd1 vssd1 vccd1 vccd1 _5570_/B sky130_fd_sc_hd__mux2_1
X_7307_ _7307_/CLK _7307_/D vssd1 vssd1 vccd1 vccd1 _7307_/Q sky130_fd_sc_hd__dfxtp_1
X_4519_ _4519_/A vssd1 vssd1 vccd1 vccd1 _7296_/D sky130_fd_sc_hd__clkbuf_1
X_7238_ _7238_/CLK _7238_/D vssd1 vssd1 vccd1 vccd1 _7238_/Q sky130_fd_sc_hd__dfxtp_1
X_5499_ _5499_/A vssd1 vssd1 vccd1 vccd1 _5499_/X sky130_fd_sc_hd__buf_1
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7169_ _7169_/CLK _7169_/D vssd1 vssd1 vccd1 vccd1 _7169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6409__526 _6410__527/A vssd1 vssd1 vccd1 vccd1 _7468_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4870_ _4828_/X _7111_/Q _4874_/S vssd1 vssd1 vccd1 vccd1 _4871_/A sky130_fd_sc_hd__mux2_1
X_3821_ _3821_/A vssd1 vssd1 vccd1 vccd1 _7590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6540_ _6535_/X _6538_/X _6539_/X vssd1 vssd1 vccd1 vccd1 _7500_/D sky130_fd_sc_hd__o21a_1
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3752_ _3752_/A vssd1 vssd1 vccd1 vccd1 _7615_/D sky130_fd_sc_hd__clkbuf_1
X_3683_ _3683_/A vssd1 vssd1 vccd1 vccd1 _7678_/D sky130_fd_sc_hd__clkbuf_1
X_6471_ _6450_/A _6159_/A _6133_/A vssd1 vssd1 vccd1 vccd1 _6474_/C sky130_fd_sc_hd__o21ai_1
XFILLER_118_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5422_ _5210_/A _5422_/B vssd1 vssd1 vccd1 vccd1 _5422_/X sky130_fd_sc_hd__and2b_1
X_5353_ _5356_/A _5352_/X _5178_/X vssd1 vssd1 vccd1 vccd1 _5353_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4304_ _4211_/X _7375_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__mux2_1
X_5284_ _5284_/A vssd1 vssd1 vccd1 vccd1 _5284_/Y sky130_fd_sc_hd__inv_2
XINSDIODE2_8 _3917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4235_ _4584_/A vssd1 vssd1 vccd1 vccd1 _4235_/X sky130_fd_sc_hd__clkbuf_4
X_7023_ _7023_/A vssd1 vssd1 vccd1 vccd1 _7728_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3082_ _6289_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3082_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4166_ _4166_/A vssd1 vssd1 vccd1 vccd1 _7428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4097_ _4119_/S vssd1 vssd1 vccd1 vccd1 _4110_/S sky130_fd_sc_hd__buf_2
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6807_ _6819_/D _6807_/B _6872_/B vssd1 vssd1 vccd1 vccd1 _6808_/A sky130_fd_sc_hd__and3b_1
X_4999_ _4999_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _5000_/A sky130_fd_sc_hd__and2_1
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6738_ _6744_/A vssd1 vssd1 vccd1 vccd1 _6738_/X sky130_fd_sc_hd__buf_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3418_ _6939_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3418_/X sky130_fd_sc_hd__clkbuf_16
X_6381__504 _6381__504/A vssd1 vssd1 vccd1 vccd1 _7446_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4020_ _4020_/A vssd1 vssd1 vccd1 vccd1 _7488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5971_ _5882_/X _5960_/X _5970_/Y vssd1 vssd1 vccd1 vccd1 _5971_/X sky130_fd_sc_hd__a21o_1
XFILLER_18_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6282__424 _6282__424/A vssd1 vssd1 vccd1 vccd1 _7366_/CLK sky130_fd_sc_hd__inv_2
X_7710_ _7710_/CLK _7710_/D vssd1 vssd1 vccd1 vccd1 _7710_/Q sky130_fd_sc_hd__dfxtp_1
X_4922_ _7051_/Q _4566_/A _4928_/S vssd1 vssd1 vccd1 vccd1 _4923_/A sky130_fd_sc_hd__mux2_1
X_7641_ _7655_/CLK _7641_/D vssd1 vssd1 vccd1 vccd1 _7641_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2720_ _5719_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2720_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4853_ _4853_/A vssd1 vssd1 vccd1 vccd1 _7119_/D sky130_fd_sc_hd__clkbuf_1
X_7572_ _7572_/CLK _7572_/D vssd1 vssd1 vccd1 vccd1 _7572_/Q sky130_fd_sc_hd__dfxtp_1
X_3804_ _7672_/Q vssd1 vssd1 vccd1 vccd1 _3804_/X sky130_fd_sc_hd__buf_6
X_4784_ _4918_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _4800_/S sky130_fd_sc_hd__nor2_2
XFILLER_118_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3735_ _3905_/A vssd1 vssd1 vccd1 vccd1 _3735_/X sky130_fd_sc_hd__buf_2
X_6523_ _6525_/A vssd1 vssd1 vccd1 vccd1 _6566_/A sky130_fd_sc_hd__buf_2
XFILLER_119_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6454_ _6454_/A _6454_/B _6454_/C _6454_/D vssd1 vssd1 vccd1 vccd1 _6455_/B sky130_fd_sc_hd__or4_1
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3666_ _3666_/A vssd1 vssd1 vccd1 vccd1 _7684_/D sky130_fd_sc_hd__clkbuf_1
X_5405_ _7532_/Q _7112_/Q _7564_/Q _7128_/Q _5303_/X _5299_/X vssd1 vssd1 vccd1 vccd1
+ _5405_/X sky130_fd_sc_hd__mux4_1
X_3597_ _7323_/Q vssd1 vssd1 vccd1 vccd1 _3597_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5336_ _5289_/A _5331_/Y _5333_/Y _5335_/Y vssd1 vssd1 vccd1 vccd1 _5337_/C sky130_fd_sc_hd__a31o_1
XFILLER_114_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5267_ _5267_/A vssd1 vssd1 vccd1 vccd1 _5365_/A sky130_fd_sc_hd__buf_2
X_4218_ _4217_/X _7406_/Q _4227_/S vssd1 vssd1 vccd1 vccd1 _4219_/A sky130_fd_sc_hd__mux2_1
X_7006_ _7006_/A vssd1 vssd1 vccd1 vccd1 _7723_/D sky130_fd_sc_hd__clkbuf_1
X_5198_ _5375_/A _7062_/Q _5376_/A input14/X vssd1 vssd1 vccd1 vccd1 _5239_/A sky130_fd_sc_hd__a22o_1
XFILLER_18_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4149_ _7435_/Q _3594_/X _4149_/S vssd1 vssd1 vccd1 vccd1 _4150_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7652_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3520_ _3520_/A vssd1 vssd1 vccd1 vccd1 _7714_/D sky130_fd_sc_hd__clkbuf_1
X_6170_ _7658_/Q _6797_/A _6170_/C _6805_/A vssd1 vssd1 vccd1 vccd1 _6171_/A sky130_fd_sc_hd__and4_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5121_ _5187_/A _5380_/B _5183_/C vssd1 vssd1 vccd1 vccd1 _5232_/B sky130_fd_sc_hd__or3_1
XFILLER_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5052_ _5052_/A vssd1 vssd1 vccd1 vccd1 _5052_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4003_ _4400_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4019_/S sky130_fd_sc_hd__nor2_4
Xclkbuf_1_0__f__2958_ clkbuf_0__2958_/X vssd1 vssd1 vccd1 vccd1 _6054__334/A sky130_fd_sc_hd__clkbuf_16
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5954_ _7539_/Q _7680_/Q _7696_/Q _7282_/Q _5907_/X _5905_/X vssd1 vssd1 vccd1 vccd1
+ _5954_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5885_ _7450_/Q _7442_/Q _7426_/Q _7418_/Q _5884_/X _4477_/A vssd1 vssd1 vccd1 vccd1
+ _5886_/B sky130_fd_sc_hd__mux4_2
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4905_ _4905_/A vssd1 vssd1 vccd1 vccd1 _7059_/D sky130_fd_sc_hd__clkbuf_1
X_7624_ _7624_/CLK _7624_/D vssd1 vssd1 vccd1 vccd1 _7624_/Q sky130_fd_sc_hd__dfxtp_1
X_4836_ _4836_/A vssd1 vssd1 vccd1 vccd1 _7125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7555_ _7555_/CLK _7555_/D vssd1 vssd1 vccd1 vccd1 _7555_/Q sky130_fd_sc_hd__dfxtp_2
X_6506_ _6482_/X _6483_/Y _6474_/X _6454_/C _6473_/Y vssd1 vssd1 vccd1 vccd1 _6509_/C
+ sky130_fd_sc_hd__a2111o_1
X_4767_ _4767_/A vssd1 vssd1 vccd1 vccd1 _7154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7486_ _7486_/CLK _7486_/D vssd1 vssd1 vccd1 vccd1 _7486_/Q sky130_fd_sc_hd__dfxtp_1
X_3718_ _3526_/X _7627_/Q _3722_/S vssd1 vssd1 vccd1 vccd1 _3719_/A sky130_fd_sc_hd__mux2_1
X_4698_ _4560_/X _7185_/Q _4706_/S vssd1 vssd1 vccd1 vccd1 _4699_/A sky130_fd_sc_hd__mux2_1
X_3649_ _3648_/X _7688_/Q _3657_/S vssd1 vssd1 vccd1 vccd1 _3650_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5319_ _5319_/A _5319_/B vssd1 vssd1 vccd1 vccd1 _5319_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6352__480 _6356__484/A vssd1 vssd1 vccd1 vccd1 _7422_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4621_ _4621_/A vssd1 vssd1 vccd1 vccd1 _7251_/D sky130_fd_sc_hd__clkbuf_1
X_6394__514 _6394__514/A vssd1 vssd1 vccd1 vccd1 _7456_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4552_ _7280_/Q _3914_/A _4552_/S vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__mux2_1
X_7340_ _7340_/CLK _7340_/D vssd1 vssd1 vccd1 vccd1 _7340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7271_ _7271_/CLK _7271_/D vssd1 vssd1 vccd1 vccd1 _7271_/Q sky130_fd_sc_hd__dfxtp_1
X_4483_ _4483_/A vssd1 vssd1 vccd1 vccd1 _6236_/C sky130_fd_sc_hd__buf_4
X_3503_ _7092_/Q _7093_/Q _7094_/Q _7091_/Q vssd1 vssd1 vccd1 vccd1 _5123_/D sky130_fd_sc_hd__or4b_1
XFILLER_89_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6222_ _6222_/A vssd1 vssd1 vccd1 vccd1 _6231_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_103_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3088_ clkbuf_0__3088_/X vssd1 vssd1 vccd1 vccd1 _6325__459/A sky130_fd_sc_hd__clkbuf_16
X_6153_ _6507_/B _6792_/D vssd1 vssd1 vccd1 vccd1 _6157_/C sky130_fd_sc_hd__xor2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _7204_/Q _5104_/B vssd1 vssd1 vccd1 vccd1 _5105_/A sky130_fd_sc_hd__and2_1
XFILLER_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5035_/A _5035_/B vssd1 vssd1 vccd1 vccd1 _5036_/A sky130_fd_sc_hd__and2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6030__314 _6030__314/A vssd1 vssd1 vccd1 vccd1 _7240_/CLK sky130_fd_sc_hd__inv_2
X_5672__232 _5674__234/A vssd1 vssd1 vccd1 vccd1 _7126_/CLK sky130_fd_sc_hd__inv_2
X_6986_ _6986_/A vssd1 vssd1 vccd1 vccd1 _7717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5937_ _5935_/X _5936_/X _5995_/S vssd1 vssd1 vccd1 vccd1 _5937_/X sky130_fd_sc_hd__mux2_2
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7607_ _7607_/CLK _7607_/D vssd1 vssd1 vccd1 vccd1 _7607_/Q sky130_fd_sc_hd__dfxtp_1
X_5868_ _6001_/A _5868_/B vssd1 vssd1 vccd1 vccd1 _5868_/X sky130_fd_sc_hd__or2_1
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4819_ _4819_/A vssd1 vssd1 vccd1 vccd1 _7130_/D sky130_fd_sc_hd__clkbuf_1
X_5799_ _5799_/A vssd1 vssd1 vccd1 vccd1 _7208_/D sky130_fd_sc_hd__clkbuf_1
X_7538_ _7538_/CLK _7538_/D vssd1 vssd1 vccd1 vccd1 _7538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7469_ _7469_/CLK _7469_/D vssd1 vssd1 vccd1 vccd1 _7469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__3294_ clkbuf_0__3294_/X vssd1 vssd1 vccd1 vccd1 _6766__17/A sky130_fd_sc_hd__clkbuf_16
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_218 vssd1 vssd1 vccd1 vccd1 CaravelHost_218/HI manufacturerID[10] sky130_fd_sc_hd__conb_1
XCaravelHost_207 vssd1 vssd1 vccd1 vccd1 CaravelHost_207/HI core1Index[7] sky130_fd_sc_hd__conb_1
XCaravelHost_229 vssd1 vssd1 vccd1 vccd1 CaravelHost_229/HI versionID[3] sky130_fd_sc_hd__conb_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5736__284 _5736__284/A vssd1 vssd1 vccd1 vccd1 _7178_/CLK sky130_fd_sc_hd__inv_2
X_6840_ _6847_/C _6843_/C vssd1 vssd1 vccd1 vccd1 _6841_/C sky130_fd_sc_hd__or2_1
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2726_ clkbuf_0__2726_/X vssd1 vssd1 vccd1 vccd1 _5803__293/A sky130_fd_sc_hd__clkbuf_16
X_6771_ _6771_/A _6771_/B vssd1 vssd1 vccd1 vccd1 _6779_/A sky130_fd_sc_hd__or2_1
XFILLER_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3983_ _4301_/C _3983_/B _3926_/A vssd1 vssd1 vccd1 vccd1 _4784_/B sky130_fd_sc_hd__or3b_4
XFILLER_31_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4604_ _4261_/X _7258_/Q _4604_/S vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__mux2_1
X_5584_ _7716_/Q _5584_/B vssd1 vssd1 vccd1 vccd1 _6234_/C sky130_fd_sc_hd__nand2_1
X_4535_ _4535_/A vssd1 vssd1 vccd1 vccd1 _7289_/D sky130_fd_sc_hd__clkbuf_1
X_7323_ _7670_/CLK _7323_/D vssd1 vssd1 vccd1 vccd1 _7323_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_104_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7254_ _7254_/CLK _7254_/D vssd1 vssd1 vccd1 vccd1 _7254_/Q sky130_fd_sc_hd__dfxtp_1
X_4466_ _3481_/X _4466_/B _4466_/C _4466_/D vssd1 vssd1 vccd1 vccd1 _4467_/C sky130_fd_sc_hd__and4b_1
X_5743__288 _5743__288/A vssd1 vssd1 vccd1 vccd1 _7182_/CLK sky130_fd_sc_hd__inv_2
X_7185_ _7185_/CLK _7185_/D vssd1 vssd1 vccd1 vccd1 _7185_/Q sky130_fd_sc_hd__dfxtp_2
X_4397_ _4395_/Y _5381_/A _4396_/X vssd1 vssd1 vccd1 vccd1 _4398_/B sky130_fd_sc_hd__o21ai_1
X_6136_ _6450_/B vssd1 vssd1 vccd1 vccd1 _6483_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5018_ _5018_/A _5024_/B vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__and2_1
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3415_ clkbuf_0__3415_/X vssd1 vssd1 vccd1 vccd1 _6930__23/A sky130_fd_sc_hd__clkbuf_16
XFILLER_60_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3277_ clkbuf_0__3277_/X vssd1 vssd1 vccd1 vccd1 _6680__123/A sky130_fd_sc_hd__clkbuf_16
XFILLER_40_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6931__24 _6931__24/A vssd1 vssd1 vccd1 vccd1 _7680_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5807__296 _5808__297/A vssd1 vssd1 vccd1 vccd1 _7214_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4320_ _7328_/Q vssd1 vssd1 vccd1 vccd1 _4320_/X sky130_fd_sc_hd__clkbuf_4
X_4251_ _4251_/A vssd1 vssd1 vccd1 vccd1 _7396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4182_ _4182_/A vssd1 vssd1 vccd1 vccd1 _7421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6211__387 _6213__389/A vssd1 vssd1 vccd1 vccd1 _7317_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__2951_ _6012_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2951_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6365__490 _6368__493/A vssd1 vssd1 vccd1 vccd1 _7432_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6765__16 _6766__17/A vssd1 vssd1 vccd1 vccd1 _7635_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6823_ _6823_/A vssd1 vssd1 vccd1 vccd1 _7643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3966_ _3981_/S vssd1 vssd1 vccd1 vccd1 _3975_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2709_ clkbuf_0__2709_/X vssd1 vssd1 vccd1 vccd1 _5668__229/A sky130_fd_sc_hd__clkbuf_16
XFILLER_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3897_ _7558_/Q _3603_/X _3897_/S vssd1 vssd1 vccd1 vccd1 _3898_/A sky130_fd_sc_hd__mux2_2
X_5636_ _5636_/A vssd1 vssd1 vccd1 vccd1 _7100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5567_ _7222_/Q _7223_/Q _7224_/Q _7225_/Q _7514_/Q _7515_/Q vssd1 vssd1 vccd1 vccd1
+ _5567_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5498_ _5498_/A vssd1 vssd1 vccd1 vccd1 _5498_/X sky130_fd_sc_hd__buf_1
X_7306_ _7306_/CLK _7306_/D vssd1 vssd1 vccd1 vccd1 _7306_/Q sky130_fd_sc_hd__dfxtp_1
X_4518_ _7296_/Q _4337_/X _4522_/S vssd1 vssd1 vccd1 vccd1 _4519_/A sky130_fd_sc_hd__mux2_1
X_7237_ _7237_/CLK _7237_/D vssd1 vssd1 vccd1 vccd1 _7237_/Q sky130_fd_sc_hd__dfxtp_1
X_4449_ _6236_/B vssd1 vssd1 vccd1 vccd1 _4486_/C sky130_fd_sc_hd__clkbuf_2
X_7168_ _7168_/CLK _7168_/D vssd1 vssd1 vccd1 vccd1 _7168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6487_/A _6119_/B _7729_/Q vssd1 vssd1 vccd1 vccd1 _6486_/B sky130_fd_sc_hd__or3_2
X_7099_ _7723_/CLK _7099_/D vssd1 vssd1 vccd1 vccd1 _7099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082__351 _6083__352/A vssd1 vssd1 vccd1 vccd1 _7280_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5685__242 _5686__243/A vssd1 vssd1 vccd1 vccd1 _7136_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3820_ _7590_/Q _3819_/X _3820_/S vssd1 vssd1 vccd1 vccd1 _3821_/A sky130_fd_sc_hd__mux2_1
X_3751_ _3750_/X _7615_/Q _3754_/S vssd1 vssd1 vccd1 vccd1 _3752_/A sky130_fd_sc_hd__mux2_1
X_3682_ _3534_/X _7678_/Q _3682_/S vssd1 vssd1 vccd1 vccd1 _3683_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6470_ _6571_/A _6777_/A _6470_/C vssd1 vssd1 vccd1 vccd1 _6470_/Y sky130_fd_sc_hd__nand3_1
X_5421_ _7121_/Q _7169_/Q _5421_/S vssd1 vssd1 vccd1 vccd1 _5422_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5352_ _7373_/Q _7344_/Q _7336_/Q _7299_/Q _4381_/A _5252_/X vssd1 vssd1 vccd1 vccd1
+ _5352_/X sky130_fd_sc_hd__mux4_2
X_4303_ _4318_/S vssd1 vssd1 vccd1 vccd1 _4312_/S sky130_fd_sc_hd__buf_2
XFILLER_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5283_ _7117_/Q _7165_/Q _5421_/S vssd1 vssd1 vccd1 vccd1 _5284_/A sky130_fd_sc_hd__mux2_1
X_7022_ _7003_/X _7022_/B vssd1 vssd1 vccd1 vccd1 _7023_/A sky130_fd_sc_hd__and2b_1
XFILLER_101_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4234_ _4234_/A vssd1 vssd1 vccd1 vccd1 _7401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3081_ _6283_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3081_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_9 _4320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4165_ _4106_/X _7428_/Q _4167_/S vssd1 vssd1 vccd1 vccd1 _4166_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _4239_/A _4175_/B vssd1 vssd1 vccd1 vccd1 _4119_/S sky130_fd_sc_hd__or2_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6806_ _6809_/A vssd1 vssd1 vccd1 vccd1 _6872_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4998_ _4998_/A vssd1 vssd1 vccd1 vccd1 _4998_/X sky130_fd_sc_hd__clkbuf_1
X_3949_ _3899_/X _7541_/Q _3957_/S vssd1 vssd1 vccd1 vccd1 _3950_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5619_ _5619_/A vssd1 vssd1 vccd1 vccd1 _7092_/D sky130_fd_sc_hd__clkbuf_1
X_6599_ _6599_/A _6599_/B _6599_/C vssd1 vssd1 vccd1 vccd1 _6600_/A sky130_fd_sc_hd__and3_1
XFILLER_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3417_ _6938_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3417_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6415__531 _6418__534/A vssd1 vssd1 vccd1 vccd1 _7473_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3279_ _6688_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3279_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6426__59 _6426__59/A vssd1 vssd1 vccd1 vccd1 _7481_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6316__451 _6319__454/A vssd1 vssd1 vccd1 vccd1 _7393_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5507__185 _5509__187/A vssd1 vssd1 vccd1 vccd1 _7041_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _5882_/A _5969_/X _5833_/X vssd1 vssd1 vccd1 vccd1 _5970_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _4921_/A vssd1 vssd1 vccd1 vccd1 _7052_/D sky130_fd_sc_hd__clkbuf_1
X_7640_ _7731_/CLK _7640_/D vssd1 vssd1 vccd1 vccd1 _7640_/Q sky130_fd_sc_hd__dfxtp_1
X_4852_ _4828_/X _7119_/Q _4856_/S vssd1 vssd1 vccd1 vccd1 _4853_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3803_ _3803_/A vssd1 vssd1 vccd1 vccd1 _7596_/D sky130_fd_sc_hd__clkbuf_1
X_7571_ _7571_/CLK _7571_/D vssd1 vssd1 vccd1 vccd1 _7571_/Q sky130_fd_sc_hd__dfxtp_1
X_4783_ _4783_/A vssd1 vssd1 vccd1 vccd1 _7146_/D sky130_fd_sc_hd__clkbuf_1
X_3734_ _3734_/A vssd1 vssd1 vccd1 vccd1 _7621_/D sky130_fd_sc_hd__clkbuf_1
X_6522_ _7498_/Q vssd1 vssd1 vccd1 vccd1 _6532_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_118_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3665_ _3664_/X _7684_/Q _3669_/S vssd1 vssd1 vccd1 vccd1 _3666_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6453_ _7501_/Q _6453_/B vssd1 vssd1 vccd1 vccd1 _6454_/D sky130_fd_sc_hd__xor2_1
XFILLER_118_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5404_ _5293_/A _5403_/X _5213_/A vssd1 vssd1 vccd1 vccd1 _5404_/X sky130_fd_sc_hd__a21o_1
X_3596_ _3596_/A vssd1 vssd1 vccd1 vccd1 _7702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5335_ _5396_/A _5334_/X _5205_/X vssd1 vssd1 vccd1 vccd1 _5335_/Y sky130_fd_sc_hd__o21ai_1
X_5266_ _5363_/A _5266_/B vssd1 vssd1 vccd1 vccd1 _5266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4217_ _4566_/A vssd1 vssd1 vccd1 vccd1 _4217_/X sky130_fd_sc_hd__buf_2
X_7005_ _7003_/X _7005_/B vssd1 vssd1 vccd1 vccd1 _7006_/A sky130_fd_sc_hd__and2b_1
X_5197_ _5450_/A vssd1 vssd1 vccd1 vccd1 _5376_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4148_ _4148_/A vssd1 vssd1 vccd1 vccd1 _7436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4079_ _4079_/A vssd1 vssd1 vccd1 vccd1 _7463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5532__201 _5532__201/A vssd1 vssd1 vccd1 vccd1 _7058_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6734__166 _6737__169/A vssd1 vssd1 vccd1 vccd1 _7610_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5730__279 _5730__279/A vssd1 vssd1 vccd1 vccd1 _7173_/CLK sky130_fd_sc_hd__inv_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5120_ _6910_/B _3511_/A vssd1 vssd1 vccd1 vccd1 _5183_/C sky130_fd_sc_hd__or2b_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5051_ _5051_/A _5057_/B vssd1 vssd1 vccd1 vccd1 _5052_/A sky130_fd_sc_hd__and2_1
XFILLER_111_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4002_ _4301_/A _4561_/B _4561_/A vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__or3b_4
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2957_ clkbuf_0__2957_/X vssd1 vssd1 vccd1 vccd1 _6046__327/A sky130_fd_sc_hd__clkbuf_16
XFILLER_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5953_ _7222_/Q _5814_/X _5952_/X _5880_/X vssd1 vssd1 vccd1 vccd1 _7222_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5884_ _5884_/A vssd1 vssd1 vccd1 vccd1 _5884_/X sky130_fd_sc_hd__buf_2
XFILLER_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4904_ _4825_/X _7059_/Q _4910_/S vssd1 vssd1 vccd1 vccd1 _4905_/A sky130_fd_sc_hd__mux2_1
X_7623_ _7623_/CLK _7623_/D vssd1 vssd1 vccd1 vccd1 _7623_/Q sky130_fd_sc_hd__dfxtp_1
X_4835_ _4834_/X _7125_/Q _4835_/S vssd1 vssd1 vccd1 vccd1 _4836_/A sky130_fd_sc_hd__mux2_1
X_7554_ _7554_/CLK _7554_/D vssd1 vssd1 vccd1 vccd1 _7554_/Q sky130_fd_sc_hd__dfxtp_2
X_4766_ _4584_/X _7154_/Q _4766_/S vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__mux2_1
X_3717_ _3717_/A vssd1 vssd1 vccd1 vccd1 _7628_/D sky130_fd_sc_hd__clkbuf_1
X_6505_ _6505_/A _6505_/B vssd1 vssd1 vccd1 vccd1 _6509_/B sky130_fd_sc_hd__or2_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7485_ _7485_/CLK _7485_/D vssd1 vssd1 vccd1 vccd1 _7485_/Q sky130_fd_sc_hd__dfxtp_1
X_4697_ _4712_/S vssd1 vssd1 vccd1 vccd1 _4706_/S sky130_fd_sc_hd__clkbuf_2
X_3648_ _4569_/A vssd1 vssd1 vccd1 vccd1 _3648_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3579_ _3927_/A _4364_/A _4385_/A vssd1 vssd1 vccd1 vccd1 _4918_/A sky130_fd_sc_hd__or3_4
XFILLER_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5318_ _7521_/Q _7158_/Q _7142_/Q _7150_/Q _4375_/A _4382_/C vssd1 vssd1 vccd1 vccd1
+ _5319_/B sky130_fd_sc_hd__mux4_1
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5249_ _7288_/Q _7074_/Q _7701_/Q _7362_/Q _5207_/X _5225_/X vssd1 vssd1 vccd1 vccd1
+ _5250_/B sky130_fd_sc_hd__mux4_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6628__81 _6628__81/A vssd1 vssd1 vccd1 vccd1 _7524_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4620_ _7251_/Q _3920_/A _4622_/S vssd1 vssd1 vccd1 vccd1 _4621_/A sky130_fd_sc_hd__mux2_1
X_4551_ _4551_/A vssd1 vssd1 vccd1 vccd1 _7281_/D sky130_fd_sc_hd__clkbuf_1
X_4482_ _4482_/A _4482_/B vssd1 vssd1 vccd1 vccd1 _7311_/D sky130_fd_sc_hd__nor2_1
X_7270_ _7270_/CLK _7270_/D vssd1 vssd1 vccd1 vccd1 _7270_/Q sky130_fd_sc_hd__dfxtp_1
X_3502_ _7104_/Q _7103_/Q vssd1 vssd1 vccd1 vccd1 _5645_/B sky130_fd_sc_hd__nor2_2
XFILLER_7_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6221_ _6221_/A vssd1 vssd1 vccd1 vccd1 _7323_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__3087_ clkbuf_0__3087_/X vssd1 vssd1 vccd1 vccd1 _6319__454/A sky130_fd_sc_hd__clkbuf_16
X_6152_ _6481_/A _7647_/Q vssd1 vssd1 vccd1 vccd1 _6792_/D sky130_fd_sc_hd__xnor2_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5103_/A vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5034_/A vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6329__461 _6331__463/A vssd1 vssd1 vccd1 vccd1 _7403_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6985_ _6981_/X _6985_/B vssd1 vssd1 vccd1 vccd1 _6986_/A sky130_fd_sc_hd__and2b_1
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5936_ _7586_/Q _7578_/Q _7570_/Q _7484_/Q _5907_/X _5908_/X vssd1 vssd1 vccd1 vccd1
+ _5936_/X sky130_fd_sc_hd__mux4_2
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7606_ _7606_/CLK _7606_/D vssd1 vssd1 vccd1 vccd1 _7606_/Q sky130_fd_sc_hd__dfxtp_2
X_5867_ _7449_/Q _7441_/Q _7425_/Q _7417_/Q _5884_/A _4462_/A vssd1 vssd1 vccd1 vccd1
+ _5868_/B sky130_fd_sc_hd__mux4_1
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4818_ _4584_/X _7130_/Q _4818_/S vssd1 vssd1 vccd1 vccd1 _4819_/A sky130_fd_sc_hd__mux2_1
X_5798_ _7208_/Q _5042_/A _5800_/S vssd1 vssd1 vccd1 vccd1 _5799_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7537_ _7537_/CLK _7537_/D vssd1 vssd1 vccd1 vccd1 _7537_/Q sky130_fd_sc_hd__dfxtp_1
X_4749_ _4749_/A vssd1 vssd1 vccd1 vccd1 _7162_/D sky130_fd_sc_hd__clkbuf_1
X_7468_ _7468_/CLK _7468_/D vssd1 vssd1 vccd1 vccd1 _7468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6419_ _6419_/A vssd1 vssd1 vccd1 vccd1 _6419_/X sky130_fd_sc_hd__buf_1
X_7399_ _7399_/CLK _7399_/D vssd1 vssd1 vccd1 vccd1 _7399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3293_ clkbuf_0__3293_/X vssd1 vssd1 vccd1 vccd1 _6761__13/A sky130_fd_sc_hd__clkbuf_16
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6943__33 _6944__34/A vssd1 vssd1 vccd1 vccd1 _7689_/CLK sky130_fd_sc_hd__inv_2
X_5649__213 _5649__213/A vssd1 vssd1 vccd1 vccd1 _7107_/CLK sky130_fd_sc_hd__inv_2
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XCaravelHost_208 vssd1 vssd1 vccd1 vccd1 CaravelHost_208/HI manufacturerID[0] sky130_fd_sc_hd__conb_1
XCaravelHost_219 vssd1 vssd1 vccd1 vccd1 CaravelHost_219/HI partID[1] sky130_fd_sc_hd__conb_1
XFILLER_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3982_ _3982_/A vssd1 vssd1 vccd1 vccd1 _7526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2725_ clkbuf_0__2725_/X vssd1 vssd1 vccd1 vccd1 _5743__288/A sky130_fd_sc_hd__clkbuf_16
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6770_ _7657_/Q _7656_/Q vssd1 vssd1 vccd1 vccd1 _6878_/B sky130_fd_sc_hd__nand2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4603_ _4603_/A vssd1 vssd1 vccd1 vccd1 _7259_/D sky130_fd_sc_hd__clkbuf_1
X_5583_ _7715_/Q vssd1 vssd1 vccd1 vccd1 _5588_/A sky130_fd_sc_hd__clkinv_2
X_4534_ _4226_/X _7289_/Q _4534_/S vssd1 vssd1 vccd1 vccd1 _4535_/A sky130_fd_sc_hd__mux2_1
X_7322_ _7670_/CLK _7322_/D vssd1 vssd1 vccd1 vccd1 _7322_/Q sky130_fd_sc_hd__dfxtp_4
X_7253_ _7253_/CLK _7253_/D vssd1 vssd1 vccd1 vccd1 _7253_/Q sky130_fd_sc_hd__dfxtp_1
X_4465_ _5884_/A vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__buf_2
X_7184_ _7184_/CLK _7184_/D vssd1 vssd1 vccd1 vccd1 _7184_/Q sky130_fd_sc_hd__dfxtp_1
X_4396_ _4396_/A vssd1 vssd1 vccd1 vccd1 _4396_/X sky130_fd_sc_hd__buf_2
X_6135_ _6149_/A _6159_/A _6135_/C vssd1 vssd1 vccd1 vccd1 _6135_/X sky130_fd_sc_hd__or3_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _5017_/A vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5919_ _7451_/Q _7443_/Q _7427_/Q _7419_/Q _5856_/X _5857_/X vssd1 vssd1 vccd1 vccd1
+ _5920_/B sky130_fd_sc_hd__mux4_1
X_6899_ _7664_/Q _6903_/B vssd1 vssd1 vccd1 vccd1 _6899_/X sky130_fd_sc_hd__or2_1
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6310__446 _6313__449/A vssd1 vssd1 vccd1 vccd1 _7388_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3276_ clkbuf_0__3276_/X vssd1 vssd1 vccd1 vccd1 _6675__119/A sky130_fd_sc_hd__clkbuf_16
XFILLER_12_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _4249_/X _7396_/Q _4253_/S vssd1 vssd1 vccd1 vccd1 _4251_/A sky130_fd_sc_hd__mux2_1
X_4181_ _4103_/X _7421_/Q _4185_/S vssd1 vssd1 vccd1 vccd1 _4182_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6822_ _6829_/C _6822_/B _6872_/B vssd1 vssd1 vccd1 vccd1 _6823_/A sky130_fd_sc_hd__and3b_1
XFILLER_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2708_ clkbuf_0__2708_/X vssd1 vssd1 vccd1 vccd1 _5661__223/A sky130_fd_sc_hd__clkbuf_16
X_3965_ _4864_/B _4846_/B vssd1 vssd1 vccd1 vccd1 _3981_/S sky130_fd_sc_hd__or2_2
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3896_ _3896_/A vssd1 vssd1 vccd1 vccd1 _7559_/D sky130_fd_sc_hd__clkbuf_1
X_5635_ _7100_/Q _7199_/Q _5635_/S vssd1 vssd1 vccd1 vccd1 _5636_/A sky130_fd_sc_hd__mux2_1
X_6179__361 _6182__364/A vssd1 vssd1 vccd1 vccd1 _7291_/CLK sky130_fd_sc_hd__inv_2
X_5566_ _7218_/Q _7219_/Q _7220_/Q _7221_/Q _7514_/Q _7515_/Q vssd1 vssd1 vccd1 vccd1
+ _5566_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5497_ _6260_/A vssd1 vssd1 vccd1 vccd1 _5497_/X sky130_fd_sc_hd__buf_1
X_7305_ _7305_/CLK _7305_/D vssd1 vssd1 vccd1 vccd1 _7305_/Q sky130_fd_sc_hd__dfxtp_1
X_4517_ _4517_/A vssd1 vssd1 vccd1 vccd1 _7297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7236_ _7236_/CLK _7236_/D vssd1 vssd1 vccd1 vccd1 _7236_/Q sky130_fd_sc_hd__dfxtp_1
X_4448_ _3671_/A _4436_/A _3822_/A vssd1 vssd1 vccd1 vccd1 _4450_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7167_ _7167_/CLK _7167_/D vssd1 vssd1 vccd1 vccd1 _7167_/Q sky130_fd_sc_hd__dfxtp_1
X_4379_ _5245_/A vssd1 vssd1 vccd1 vccd1 _5421_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_86_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6118_ _6118_/A vssd1 vssd1 vccd1 vccd1 _6816_/A sky130_fd_sc_hd__clkbuf_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7727_/CLK _7098_/D vssd1 vssd1 vccd1 vccd1 _7098_/Q sky130_fd_sc_hd__dfxtp_1
X_6049_ _6049_/A vssd1 vssd1 vccd1 vccd1 _6049_/X sky130_fd_sc_hd__buf_1
XFILLER_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5500__180 _5502__182/A vssd1 vssd1 vccd1 vccd1 _7036_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3750_ _3920_/A vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__buf_2
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3681_ _3681_/A vssd1 vssd1 vccd1 vccd1 _7679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5420_ _5131_/X _5413_/X _5415_/X _5419_/X _5161_/A vssd1 vssd1 vccd1 vccd1 _5420_/X
+ sky130_fd_sc_hd__a311o_1
X_5351_ _5351_/A _5351_/B vssd1 vssd1 vccd1 vccd1 _5351_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5282_ _5365_/A vssd1 vssd1 vccd1 vccd1 _5291_/A sky130_fd_sc_hd__clkbuf_2
X_4302_ _4802_/A _4506_/B vssd1 vssd1 vccd1 vccd1 _4318_/S sky130_fd_sc_hd__or2_2
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4233_ _4232_/X _7401_/Q _4236_/S vssd1 vssd1 vccd1 vccd1 _4234_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7021_ _6917_/A _6784_/A _7024_/S vssd1 vssd1 vccd1 vccd1 _7022_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3080_ _6277_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3080_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4164_ _4164_/A vssd1 vssd1 vccd1 vccd1 _7429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4095_ _4095_/A _4095_/B _3900_/C vssd1 vssd1 vccd1 vccd1 _4175_/B sky130_fd_sc_hd__or3b_1
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6805_ _6805_/A _6864_/A vssd1 vssd1 vccd1 vccd1 _6809_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4997_ _4997_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _4998_/A sky130_fd_sc_hd__and2_1
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3948_ _3963_/S vssd1 vssd1 vccd1 vccd1 _3957_/S sky130_fd_sc_hd__clkbuf_2
X_3879_ _3879_/A vssd1 vssd1 vccd1 vccd1 _7566_/D sky130_fd_sc_hd__clkbuf_1
X_5618_ _7092_/Q _5075_/A _5624_/S vssd1 vssd1 vccd1 vccd1 _5619_/A sky130_fd_sc_hd__mux2_1
X_6598_ _6561_/A _6498_/A _6597_/Y _6534_/A vssd1 vssd1 vccd1 vccd1 _6599_/C sky130_fd_sc_hd__a22o_1
XFILLER_117_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3416_ _6932_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3416_/X sky130_fd_sc_hd__clkbuf_16
X_5549_ _5549_/A vssd1 vssd1 vccd1 vccd1 _7066_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3278_ _6682_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3278_/X sky130_fd_sc_hd__clkbuf_16
X_7219_ _7516_/CLK _7219_/D vssd1 vssd1 vccd1 vccd1 _7219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2630_ clkbuf_0__2630_/X vssd1 vssd1 vccd1 vccd1 _5509__187/A sky130_fd_sc_hd__clkbuf_16
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4920_ _7052_/Q _4560_/A _4928_/S vssd1 vssd1 vccd1 vccd1 _4921_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4851_ _4851_/A vssd1 vssd1 vccd1 vccd1 _7120_/D sky130_fd_sc_hd__clkbuf_1
X_3802_ _7596_/Q _3801_/X _3811_/S vssd1 vssd1 vccd1 vccd1 _3803_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7570_ _7570_/CLK _7570_/D vssd1 vssd1 vccd1 vccd1 _7570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4782_ _7146_/Q _4343_/X _4782_/S vssd1 vssd1 vccd1 vccd1 _4783_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3733_ _3730_/X _7621_/Q _3745_/S vssd1 vssd1 vccd1 vccd1 _3734_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6521_ _6579_/B _6579_/C _6520_/Y _5991_/X vssd1 vssd1 vccd1 vccd1 _7497_/D sky130_fd_sc_hd__o211a_1
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3664_ _4581_/A vssd1 vssd1 vccd1 vccd1 _3664_/X sky130_fd_sc_hd__buf_2
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6452_ _6452_/A _6452_/B vssd1 vssd1 vccd1 vccd1 _6453_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5403_ _7689_/Q _7612_/Q _5403_/S vssd1 vssd1 vccd1 vccd1 _5403_/X sky130_fd_sc_hd__mux2_1
X_3595_ _7702_/Q _3594_/X _3595_/S vssd1 vssd1 vccd1 vccd1 _3596_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5334_ _7134_/Q _7057_/Q _7049_/Q _7270_/Q _5303_/X _5299_/X vssd1 vssd1 vccd1 vccd1
+ _5334_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5265_ _7156_/Q _7148_/Q _5362_/S vssd1 vssd1 vccd1 vccd1 _5266_/B sky130_fd_sc_hd__mux2_1
X_4216_ _4216_/A vssd1 vssd1 vccd1 vccd1 _7407_/D sky130_fd_sc_hd__clkbuf_1
X_5196_ _5458_/A vssd1 vssd1 vccd1 vccd1 _5375_/A sky130_fd_sc_hd__clkbuf_4
X_7004_ _4995_/A _6137_/A _7007_/S vssd1 vssd1 vccd1 vccd1 _7005_/B sky130_fd_sc_hd__mux2_1
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4147_ _7436_/Q _3591_/X _4149_/S vssd1 vssd1 vccd1 vccd1 _4148_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4078_ _7463_/Q _3794_/X _4086_/S vssd1 vssd1 vccd1 vccd1 _4079_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6431__63 _6432__64/A vssd1 vssd1 vccd1 vccd1 _7485_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6719_ _6719_/A vssd1 vssd1 vccd1 vccd1 _6719_/X sky130_fd_sc_hd__buf_1
X_7699_ _7699_/CLK _7699_/D vssd1 vssd1 vccd1 vccd1 _7699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _5050_/A vssd1 vssd1 vccd1 vccd1 _5050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5698__253 _5698__253/A vssd1 vssd1 vccd1 vccd1 _7147_/CLK sky130_fd_sc_hd__inv_2
X_4001_ _4001_/A vssd1 vssd1 vccd1 vccd1 _7517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2956_ clkbuf_0__2956_/X vssd1 vssd1 vccd1 vccd1 _6042__324/A sky130_fd_sc_hd__clkbuf_16
XFILLER_65_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5952_ _5882_/X _5941_/X _5951_/Y vssd1 vssd1 vccd1 vccd1 _5952_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4903_ _4903_/A vssd1 vssd1 vccd1 vccd1 _7060_/D sky130_fd_sc_hd__clkbuf_1
X_5883_ _5910_/A vssd1 vssd1 vccd1 vccd1 _5966_/A sky130_fd_sc_hd__clkbuf_2
X_7622_ _7622_/CLK _7622_/D vssd1 vssd1 vccd1 vccd1 _7622_/Q sky130_fd_sc_hd__dfxtp_1
X_4834_ _7324_/Q vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__buf_2
X_7553_ _7553_/CLK _7553_/D vssd1 vssd1 vccd1 vccd1 _7553_/Q sky130_fd_sc_hd__dfxtp_1
X_4765_ _4765_/A vssd1 vssd1 vccd1 vccd1 _7155_/D sky130_fd_sc_hd__clkbuf_1
X_3716_ _3522_/X _7628_/Q _3722_/S vssd1 vssd1 vccd1 vccd1 _3717_/A sky130_fd_sc_hd__mux2_1
X_6504_ _6504_/A _6504_/B _6504_/C _6504_/D vssd1 vssd1 vccd1 vccd1 _6504_/X sky130_fd_sc_hd__or4_1
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7484_ _7484_/CLK _7484_/D vssd1 vssd1 vccd1 vccd1 _7484_/Q sky130_fd_sc_hd__dfxtp_1
X_4696_ _4821_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4712_/S sky130_fd_sc_hd__or2_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _7326_/Q vssd1 vssd1 vccd1 vccd1 _4569_/A sky130_fd_sc_hd__clkbuf_4
X_3578_ _6913_/A _3513_/A _3611_/A vssd1 vssd1 vccd1 vccd1 _4385_/A sky130_fd_sc_hd__a21o_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5317_ _5319_/A _5317_/B vssd1 vssd1 vccd1 vccd1 _5317_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5248_ _5244_/X _5246_/X _5349_/S vssd1 vssd1 vccd1 vccd1 _5248_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5179_ _5289_/A _5172_/X _5177_/X _5178_/X vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__o211a_1
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6740__171 _6743__174/A vssd1 vssd1 vccd1 vccd1 _7615_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4550_ _7281_/Q _3911_/A _4552_/S vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__mux2_1
X_4481_ _4477_/A _4477_/B _4438_/X vssd1 vssd1 vccd1 vccd1 _4482_/B sky130_fd_sc_hd__o21ai_1
XFILLER_7_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3501_ _7083_/Q _7084_/Q _7089_/Q _7090_/Q vssd1 vssd1 vccd1 vccd1 _3501_/X sky130_fd_sc_hd__or4_4
XFILLER_116_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6220_ _7661_/Q _6220_/B vssd1 vssd1 vccd1 vccd1 _6221_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_0__f__3086_ clkbuf_0__3086_/X vssd1 vssd1 vccd1 vccd1 _6312__448/A sky130_fd_sc_hd__clkbuf_16
X_6151_ _6151_/A vssd1 vssd1 vccd1 vccd1 _6507_/B sky130_fd_sc_hd__buf_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5102_ _5555_/B _7203_/Q _5102_/C _5102_/D vssd1 vssd1 vccd1 vccd1 _5103_/A sky130_fd_sc_hd__and4_4
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6683__125 _6685__127/A vssd1 vssd1 vccd1 vccd1 _7569_/CLK sky130_fd_sc_hd__inv_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A _5035_/B vssd1 vssd1 vccd1 vccd1 _5034_/A sky130_fd_sc_hd__and2_1
XFILLER_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6634__85 _6637__88/A vssd1 vssd1 vccd1 vccd1 _7529_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6984_ _5008_/A _6463_/A _7000_/S vssd1 vssd1 vccd1 vccd1 _6985_/B sky130_fd_sc_hd__mux2_1
X_5935_ _7538_/Q _7679_/Q _7695_/Q _7281_/Q _5851_/X _5905_/X vssd1 vssd1 vccd1 vccd1
+ _5935_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5866_ _5910_/A vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__clkbuf_2
X_7605_ _7605_/CLK _7605_/D vssd1 vssd1 vccd1 vccd1 _7605_/Q sky130_fd_sc_hd__dfxtp_1
X_4817_ _4817_/A vssd1 vssd1 vccd1 vccd1 _7131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5797_ _5797_/A vssd1 vssd1 vccd1 vccd1 _7207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7536_ _7536_/CLK _7536_/D vssd1 vssd1 vccd1 vccd1 _7536_/Q sky130_fd_sc_hd__dfxtp_1
X_4748_ _7162_/Q _4343_/X _4748_/S vssd1 vssd1 vccd1 vccd1 _4749_/A sky130_fd_sc_hd__mux2_1
X_7467_ _7467_/CLK _7467_/D vssd1 vssd1 vccd1 vccd1 _7467_/Q sky130_fd_sc_hd__dfxtp_1
X_4679_ _4694_/S vssd1 vssd1 vccd1 vccd1 _4688_/S sky130_fd_sc_hd__clkbuf_4
X_7398_ _7398_/CLK _7398_/D vssd1 vssd1 vccd1 vccd1 _7398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__3292_ clkbuf_0__3292_/X vssd1 vssd1 vccd1 vccd1 _6754__7/A sky130_fd_sc_hd__clkbuf_16
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_209 vssd1 vssd1 vccd1 vccd1 CaravelHost_209/HI manufacturerID[1] sky130_fd_sc_hd__conb_1
XFILLER_106_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6747__177 _6747__177/A vssd1 vssd1 vccd1 vccd1 _7621_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__2724_ clkbuf_0__2724_/X vssd1 vssd1 vccd1 vccd1 _5745_/A sky130_fd_sc_hd__clkbuf_16
X_3981_ _3668_/X _7526_/Q _3981_/S vssd1 vssd1 vccd1 vccd1 _3982_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5651_ _5669_/A vssd1 vssd1 vccd1 vccd1 _5651_/X sky130_fd_sc_hd__buf_1
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4602_ _4258_/X _7259_/Q _4604_/S vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4533_ _4533_/A vssd1 vssd1 vccd1 vccd1 _7290_/D sky130_fd_sc_hd__clkbuf_1
X_7321_ _7670_/CLK _7321_/D vssd1 vssd1 vccd1 vccd1 _7321_/Q sky130_fd_sc_hd__dfxtp_4
X_7252_ _7252_/CLK _7252_/D vssd1 vssd1 vccd1 vccd1 _7252_/Q sky130_fd_sc_hd__dfxtp_1
X_4464_ _5856_/A vssd1 vssd1 vccd1 vccd1 _5884_/A sky130_fd_sc_hd__buf_4
X_7183_ _7183_/CLK _7183_/D vssd1 vssd1 vccd1 vccd1 _7183_/Q sky130_fd_sc_hd__dfxtp_1
X_4395_ _7359_/Q vssd1 vssd1 vccd1 vccd1 _4395_/Y sky130_fd_sc_hd__inv_2
X_6134_ _6450_/A _6452_/A _6135_/C vssd1 vssd1 vccd1 vccd1 _6134_/Y sky130_fd_sc_hd__o21ai_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5016_/A _5024_/B vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__and2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6069__345 _6079__349/A vssd1 vssd1 vccd1 vccd1 _7271_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6622__77 _6624__79/A vssd1 vssd1 vccd1 vccd1 _7520_/CLK sky130_fd_sc_hd__inv_2
X_5918_ _5911_/X _5916_/X _5999_/S vssd1 vssd1 vccd1 vccd1 _5918_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6898_ _7663_/Q _6892_/X _6897_/X _6880_/X vssd1 vssd1 vccd1 vccd1 _7662_/D sky130_fd_sc_hd__o211a_1
XFILLER_42_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6377__500 _6379__502/A vssd1 vssd1 vccd1 vccd1 _7442_/CLK sky130_fd_sc_hd__inv_2
X_5849_ _7218_/Q _5814_/X _5848_/X vssd1 vssd1 vccd1 vccd1 _7218_/D sky130_fd_sc_hd__o21ba_1
XFILLER_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7519_ _7519_/CLK _7519_/D vssd1 vssd1 vccd1 vccd1 _7519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6013__300 _6015__302/A vssd1 vssd1 vccd1 vccd1 _7226_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3275_ clkbuf_0__3275_/X vssd1 vssd1 vccd1 vccd1 _6666__111/A sky130_fd_sc_hd__clkbuf_16
X_6278__420 _6282__424/A vssd1 vssd1 vccd1 vccd1 _7362_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4180_ _4180_/A vssd1 vssd1 vccd1 vccd1 _7422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6821_ _6821_/A _6821_/B vssd1 vssd1 vccd1 vccd1 _6822_/B sky130_fd_sc_hd__or2_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2707_ clkbuf_0__2707_/X vssd1 vssd1 vccd1 vccd1 _5656__219/A sky130_fd_sc_hd__clkbuf_16
X_3964_ _3964_/A vssd1 vssd1 vccd1 vccd1 _7534_/D sky130_fd_sc_hd__clkbuf_1
X_3895_ _7559_/Q _3600_/X _3897_/S vssd1 vssd1 vccd1 vccd1 _3896_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__2638_ clkbuf_0__2638_/X vssd1 vssd1 vccd1 vccd1 _5572__204/A sky130_fd_sc_hd__clkbuf_16
X_5634_ _5634_/A vssd1 vssd1 vccd1 vccd1 _7099_/D sky130_fd_sc_hd__clkbuf_1
X_7304_ _7304_/CLK _7304_/D vssd1 vssd1 vccd1 vccd1 _7304_/Q sky130_fd_sc_hd__dfxtp_1
X_5565_ _6599_/A vssd1 vssd1 vccd1 vccd1 _6569_/A sky130_fd_sc_hd__buf_2
XFILLER_117_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5496_ _5496_/A vssd1 vssd1 vccd1 vccd1 _5496_/X sky130_fd_sc_hd__buf_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4516_ _7297_/Q _4334_/X _4516_/S vssd1 vssd1 vccd1 vccd1 _4517_/A sky130_fd_sc_hd__mux2_1
X_7235_ _7235_/CLK _7235_/D vssd1 vssd1 vccd1 vccd1 _7235_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3294_ _6763_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3294_/X sky130_fd_sc_hd__clkbuf_16
X_4447_ _4447_/A _4447_/B vssd1 vssd1 vccd1 vccd1 _7317_/D sky130_fd_sc_hd__nor2_1
X_6372__496 _6373__497/A vssd1 vssd1 vccd1 vccd1 _7438_/CLK sky130_fd_sc_hd__inv_2
X_7166_ _7166_/CLK _7166_/D vssd1 vssd1 vccd1 vccd1 _7166_/Q sky130_fd_sc_hd__dfxtp_1
X_6117_ _7642_/Q vssd1 vssd1 vccd1 vccd1 _6118_/A sky130_fd_sc_hd__inv_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4378_ _7347_/Q vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6438__69 _6438__69/A vssd1 vssd1 vccd1 vccd1 _7491_/CLK sky130_fd_sc_hd__inv_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7723_/CLK _7097_/D vssd1 vssd1 vccd1 vccd1 _7097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6696__135 _6700__139/A vssd1 vssd1 vccd1 vccd1 _7579_/CLK sky130_fd_sc_hd__inv_2
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7731_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5692__248 _5693__249/A vssd1 vssd1 vccd1 vccd1 _7142_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3680_ _3530_/X _7679_/Q _3682_/S vssd1 vssd1 vccd1 vccd1 _3681_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5350_ _7291_/Q _7077_/Q _7704_/Q _7365_/Q _5207_/X _5225_/X vssd1 vssd1 vccd1 vccd1
+ _5351_/B sky130_fd_sc_hd__mux4_1
XFILLER_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5281_ _7729_/Q vssd1 vssd1 vccd1 vccd1 _5281_/X sky130_fd_sc_hd__clkbuf_4
X_4301_ _4301_/A _4561_/A _4301_/C vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__nand3_4
X_4232_ _4581_/A vssd1 vssd1 vccd1 vccd1 _4232_/X sky130_fd_sc_hd__buf_2
X_7020_ _7020_/A vssd1 vssd1 vccd1 vccd1 _7727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4163_ _4103_/X _7429_/Q _4167_/S vssd1 vssd1 vccd1 vccd1 _4164_/A sky130_fd_sc_hd__mux2_1
X_4094_ _7674_/Q vssd1 vssd1 vccd1 vccd1 _4094_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4996_ _4996_/A vssd1 vssd1 vccd1 vccd1 _4996_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6804_ _6803_/B _6794_/B _6797_/A vssd1 vssd1 vccd1 vccd1 _6864_/A sky130_fd_sc_hd__a21bo_1
X_3947_ _4542_/B _4678_/A vssd1 vssd1 vccd1 vccd1 _3963_/S sky130_fd_sc_hd__nand2_4
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3878_ _3753_/X _7566_/Q _3878_/S vssd1 vssd1 vccd1 vccd1 _3879_/A sky130_fd_sc_hd__mux2_1
X_5617_ _5617_/A vssd1 vssd1 vccd1 vccd1 _7091_/D sky130_fd_sc_hd__clkbuf_1
X_6597_ _7511_/Q _6604_/C vssd1 vssd1 vccd1 vccd1 _6597_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_0__3415_ _6926_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3415_/X sky130_fd_sc_hd__clkbuf_16
X_5548_ _6919_/A _7066_/Q _5552_/S vssd1 vssd1 vccd1 vccd1 _5549_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7218_ _7516_/CLK _7218_/D vssd1 vssd1 vccd1 vccd1 _7218_/Q sky130_fd_sc_hd__dfxtp_1
X_5479_ _5474_/X _7199_/Q input16/X _5475_/X vssd1 vssd1 vccd1 vccd1 _5479_/X sky130_fd_sc_hd__a22o_2
Xclkbuf_0__3277_ _6676_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3277_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7149_ _7149_/CLK _7149_/D vssd1 vssd1 vccd1 vccd1 _7149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6704__142 _6704__142/A vssd1 vssd1 vccd1 vccd1 _7586_/CLK sky130_fd_sc_hd__inv_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3112_ clkbuf_0__3112_/X vssd1 vssd1 vccd1 vccd1 _6441__71/A sky130_fd_sc_hd__clkbuf_16
XFILLER_80_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6240__393 _6240__393/A vssd1 vssd1 vccd1 vccd1 _7333_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _4825_/X _7120_/Q _4856_/S vssd1 vssd1 vccd1 vccd1 _4851_/A sky130_fd_sc_hd__mux2_1
X_6026__310 _6027__311/A vssd1 vssd1 vccd1 vccd1 _7236_/CLK sky130_fd_sc_hd__inv_2
X_3801_ _7673_/Q vssd1 vssd1 vccd1 vccd1 _3801_/X sky130_fd_sc_hd__buf_6
X_6323__457 _6323__457/A vssd1 vssd1 vccd1 vccd1 _7399_/CLK sky130_fd_sc_hd__inv_2
X_4781_ _4781_/A vssd1 vssd1 vccd1 vccd1 _7147_/D sky130_fd_sc_hd__clkbuf_1
X_6520_ _6579_/B _6579_/C vssd1 vssd1 vccd1 vccd1 _6520_/Y sky130_fd_sc_hd__nand2_1
X_3732_ _3754_/S vssd1 vssd1 vccd1 vccd1 _3745_/S sky130_fd_sc_hd__buf_2
XFILLER_119_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3663_ _7322_/Q vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__buf_2
X_6451_ _7502_/Q _6451_/B vssd1 vssd1 vccd1 vccd1 _6454_/C sky130_fd_sc_hd__xnor2_1
X_6382_ _6382_/A vssd1 vssd1 vccd1 vccd1 _6382_/X sky130_fd_sc_hd__buf_1
X_5402_ _4396_/A _7168_/Q _5401_/X vssd1 vssd1 vccd1 vccd1 _5402_/X sky130_fd_sc_hd__o21a_1
X_5333_ _7436_/Q _4396_/X _5332_/X vssd1 vssd1 vccd1 vccd1 _5333_/Y sky130_fd_sc_hd__o21ai_1
X_3594_ _7324_/Q vssd1 vssd1 vccd1 vccd1 _3594_/X sky130_fd_sc_hd__buf_4
X_5264_ _5418_/A vssd1 vssd1 vccd1 vccd1 _5264_/X sky130_fd_sc_hd__buf_2
XFILLER_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4215_ _4211_/X _7407_/Q _4227_/S vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__mux2_1
X_5195_ _5112_/X _5190_/X _5194_/X vssd1 vssd1 vccd1 vccd1 _5195_/X sky130_fd_sc_hd__a21o_1
X_7003_ _7034_/A vssd1 vssd1 vccd1 vccd1 _7003_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4146_ _4146_/A vssd1 vssd1 vccd1 vccd1 _7437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4092_/S vssd1 vssd1 vccd1 vccd1 _4086_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4979_ _6913_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4980_/A sky130_fd_sc_hd__and2_1
XFILLER_51_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7698_ _7698_/CLK _7698_/D vssd1 vssd1 vccd1 vccd1 _7698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4000_ _3668_/X _7517_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _4001_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2955_ clkbuf_0__2955_/X vssd1 vssd1 vccd1 vccd1 _6035__318/A sky130_fd_sc_hd__clkbuf_16
XFILLER_53_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5951_ _5902_/A _5950_/X _5833_/X vssd1 vssd1 vccd1 vccd1 _5951_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4902_ _4820_/X _7060_/Q _4910_/S vssd1 vssd1 vccd1 vccd1 _4903_/A sky130_fd_sc_hd__mux2_1
X_5882_ _5882_/A vssd1 vssd1 vccd1 vccd1 _5882_/X sky130_fd_sc_hd__clkbuf_2
X_6247__399 _6247__399/A vssd1 vssd1 vccd1 vccd1 _7339_/CLK sky130_fd_sc_hd__inv_2
X_7621_ _7621_/CLK _7621_/D vssd1 vssd1 vccd1 vccd1 _7621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4833_ _4833_/A vssd1 vssd1 vccd1 vccd1 _7126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7552_ _7552_/CLK _7552_/D vssd1 vssd1 vccd1 vccd1 _7552_/Q sky130_fd_sc_hd__dfxtp_1
X_4764_ _4581_/X _7155_/Q _4766_/S vssd1 vssd1 vccd1 vccd1 _4765_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7483_ _7483_/CLK _7483_/D vssd1 vssd1 vccd1 vccd1 _7483_/Q sky130_fd_sc_hd__dfxtp_1
X_3715_ _3715_/A vssd1 vssd1 vccd1 vccd1 _7629_/D sky130_fd_sc_hd__clkbuf_1
X_6503_ _7510_/Q _6503_/B vssd1 vssd1 vccd1 vccd1 _6504_/C sky130_fd_sc_hd__xnor2_1
XFILLER_119_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4695_ _4695_/A vssd1 vssd1 vccd1 vccd1 _7210_/D sky130_fd_sc_hd__clkbuf_1
X_3646_ _3646_/A vssd1 vssd1 vccd1 vccd1 _7689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3577_ _3577_/A vssd1 vssd1 vccd1 vccd1 _6913_/A sky130_fd_sc_hd__buf_8
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6296_ _6320_/A vssd1 vssd1 vccd1 vccd1 _6296_/X sky130_fd_sc_hd__buf_1
X_5316_ _7118_/Q _7166_/Q _7687_/Q _7610_/Q _5171_/X _5291_/A vssd1 vssd1 vccd1 vccd1
+ _5317_/B sky130_fd_sc_hd__mux4_1
X_5247_ _5262_/A vssd1 vssd1 vccd1 vccd1 _5349_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5178_ _5178_/A vssd1 vssd1 vccd1 vccd1 _5178_/X sky130_fd_sc_hd__clkbuf_2
X_4129_ _4106_/X _7444_/Q _4131_/S vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6955__43 _6955__43/A vssd1 vssd1 vccd1 vccd1 _7699_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3500_ _3511_/A _6910_/B vssd1 vssd1 vccd1 vccd1 _5185_/B sky130_fd_sc_hd__or2_2
X_4480_ _4480_/A vssd1 vssd1 vccd1 vccd1 _7312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3085_ clkbuf_0__3085_/X vssd1 vssd1 vccd1 vccd1 _6307__444/A sky130_fd_sc_hd__clkbuf_16
X_6150_ _7725_/Q _6446_/A _6483_/C vssd1 vssd1 vccd1 vccd1 _6151_/A sky130_fd_sc_hd__or3b_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6173__357 _6173__357/A vssd1 vssd1 vccd1 vccd1 _7287_/CLK sky130_fd_sc_hd__inv_2
X_5101_ _5450_/A vssd1 vssd1 vccd1 vccd1 _5102_/D sky130_fd_sc_hd__buf_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_10_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7655_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5032_/A vssd1 vssd1 vccd1 vccd1 _5032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6983_ _7007_/S vssd1 vssd1 vccd1 vccd1 _7000_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_25_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5934_ _7221_/Q _5814_/X _5933_/X _5880_/X vssd1 vssd1 vccd1 vccd1 _7221_/D sky130_fd_sc_hd__o211a_1
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5865_ _5854_/X _5859_/X _5864_/X _4473_/A _5832_/A vssd1 vssd1 vccd1 vccd1 _5865_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7604_ _7604_/CLK _7604_/D vssd1 vssd1 vccd1 vccd1 _7604_/Q sky130_fd_sc_hd__dfxtp_2
X_4816_ _4581_/X _7131_/Q _4818_/S vssd1 vssd1 vccd1 vccd1 _4817_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5796_ _7207_/Q _5040_/A _5800_/S vssd1 vssd1 vccd1 vccd1 _5797_/A sky130_fd_sc_hd__mux2_1
X_7535_ _7535_/CLK _7535_/D vssd1 vssd1 vccd1 vccd1 _7535_/Q sky130_fd_sc_hd__dfxtp_1
X_4747_ _4747_/A vssd1 vssd1 vccd1 vccd1 _7163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7466_ _7466_/CLK _7466_/D vssd1 vssd1 vccd1 vccd1 _7466_/Q sky130_fd_sc_hd__dfxtp_1
X_4678_ _4678_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4694_/S sky130_fd_sc_hd__nand2_2
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3629_ _3629_/A vssd1 vssd1 vccd1 vccd1 _7692_/D sky130_fd_sc_hd__clkbuf_1
X_7397_ _7397_/CLK _7397_/D vssd1 vssd1 vccd1 vccd1 _7397_/Q sky130_fd_sc_hd__dfxtp_1
X_6336__467 _6338__469/A vssd1 vssd1 vccd1 vccd1 _7409_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6928__21 _6931__24/A vssd1 vssd1 vccd1 vccd1 _7677_/CLK sky130_fd_sc_hd__inv_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__3291_ clkbuf_0__3291_/X vssd1 vssd1 vccd1 vccd1 _6763_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_72_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5656__219 _5656__219/A vssd1 vssd1 vccd1 vccd1 _7113_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3980_ _3980_/A vssd1 vssd1 vccd1 vccd1 _7527_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__2723_ clkbuf_0__2723_/X vssd1 vssd1 vccd1 vccd1 _6207_/A sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4601_ _4601_/A vssd1 vssd1 vccd1 vccd1 _7260_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4532_ _4223_/X _7290_/Q _4534_/S vssd1 vssd1 vccd1 vccd1 _4533_/A sky130_fd_sc_hd__mux2_1
X_7320_ _7320_/CLK _7320_/D vssd1 vssd1 vccd1 vccd1 _7320_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7251_ _7251_/CLK _7251_/D vssd1 vssd1 vccd1 vccd1 _7251_/Q sky130_fd_sc_hd__dfxtp_1
X_4463_ _7310_/Q vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7182_ _7182_/CLK _7182_/D vssd1 vssd1 vccd1 vccd1 _7182_/Q sky130_fd_sc_hd__dfxtp_1
X_4394_ _6274_/A _4394_/B _4394_/C vssd1 vssd1 vccd1 vccd1 _7348_/D sky130_fd_sc_hd__nor3_1
X_6133_ _6133_/A _7645_/Q vssd1 vssd1 vccd1 vccd1 _6135_/C sky130_fd_sc_hd__xnor2_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5015_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5024_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5917_ _5917_/A vssd1 vssd1 vccd1 vccd1 _5999_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6897_ _7662_/Q _6905_/B vssd1 vssd1 vccd1 vccd1 _6897_/X sky130_fd_sc_hd__or2_1
XFILLER_34_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5848_ _5832_/Y _5833_/X _5846_/Y _6607_/A vssd1 vssd1 vccd1 vccd1 _5848_/X sky130_fd_sc_hd__a31o_1
X_5779_ _5779_/A vssd1 vssd1 vccd1 vccd1 _7199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7518_ _7518_/CLK _7518_/D vssd1 vssd1 vccd1 vccd1 _7518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7449_ _7449_/CLK _7449_/D vssd1 vssd1 vccd1 vccd1 _7449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5575__206 _5576__207/A vssd1 vssd1 vccd1 vccd1 _7074_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__3274_ clkbuf_0__3274_/X vssd1 vssd1 vccd1 vccd1 _6663__109/A sky130_fd_sc_hd__clkbuf_16
XFILLER_9_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6820_ _6833_/D vssd1 vssd1 vccd1 vccd1 _6829_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3963_ _3923_/X _7534_/Q _3963_/S vssd1 vssd1 vccd1 vccd1 _3964_/A sky130_fd_sc_hd__mux2_1
X_6751_ _6763_/A vssd1 vssd1 vccd1 vccd1 _6751_/X sky130_fd_sc_hd__buf_1
X_5517__189 _5517__189/A vssd1 vssd1 vccd1 vccd1 _7046_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6682_ _6682_/A vssd1 vssd1 vccd1 vccd1 _6682_/X sky130_fd_sc_hd__buf_1
X_3894_ _3894_/A vssd1 vssd1 vccd1 vccd1 _7560_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__2637_ clkbuf_0__2637_/X vssd1 vssd1 vccd1 vccd1 _5529__199/A sky130_fd_sc_hd__clkbuf_16
X_5633_ _7099_/Q _7198_/Q _5635_/S vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5564_ _6911_/A _3513_/X _6993_/A vssd1 vssd1 vccd1 vccd1 _6599_/A sky130_fd_sc_hd__a21oi_4
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7303_ _7303_/CLK _7303_/D vssd1 vssd1 vccd1 vccd1 _7303_/Q sky130_fd_sc_hd__dfxtp_1
X_4515_ _4515_/A vssd1 vssd1 vccd1 vccd1 _7298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5495_ _5495_/A vssd1 vssd1 vccd1 vccd1 _5495_/X sky130_fd_sc_hd__clkbuf_1
X_7234_ _7234_/CLK _7234_/D vssd1 vssd1 vccd1 vccd1 _7234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3293_ _6757_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3293_/X sky130_fd_sc_hd__clkbuf_16
X_4446_ _4039_/C _4606_/B _4438_/X vssd1 vssd1 vccd1 vccd1 _4447_/B sky130_fd_sc_hd__o21ai_1
X_7165_ _7165_/CLK _7165_/D vssd1 vssd1 vccd1 vccd1 _7165_/Q sky130_fd_sc_hd__dfxtp_1
X_4377_ _5230_/A _4377_/B vssd1 vssd1 vccd1 vccd1 _5381_/A sky130_fd_sc_hd__and2_2
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6116_ _6100_/Y _6101_/X _6778_/B _6778_/A _6771_/A vssd1 vssd1 vccd1 vccd1 _6165_/A
+ sky130_fd_sc_hd__a2111o_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7723_/CLK _7096_/D vssd1 vssd1 vccd1 vccd1 _7096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6186__367 _6186__367/A vssd1 vssd1 vccd1 vccd1 _7297_/CLK sky130_fd_sc_hd__inv_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5726__275 _5728__277/A vssd1 vssd1 vccd1 vccd1 _7169_/CLK sky130_fd_sc_hd__inv_2
X_5581__210 _5649__213/A vssd1 vssd1 vccd1 vccd1 _7078_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5280_ _5375_/A _7064_/Q _5376_/A input28/X vssd1 vssd1 vccd1 vccd1 _5311_/A sky130_fd_sc_hd__a22o_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4300_ _4300_/A vssd1 vssd1 vccd1 vccd1 _7376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4231_ _4231_/A vssd1 vssd1 vccd1 vccd1 _7402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4162_ _4162_/A vssd1 vssd1 vccd1 vccd1 _7430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4093_ _4093_/A vssd1 vssd1 vccd1 vccd1 _7456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6443__73 _6618__74/A vssd1 vssd1 vccd1 vccd1 _7495_/CLK sky130_fd_sc_hd__inv_2
X_4995_ _4995_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _4996_/A sky130_fd_sc_hd__and2_1
X_6803_ _7640_/Q _6803_/B _6781_/A vssd1 vssd1 vccd1 vccd1 _6807_/B sky130_fd_sc_hd__or3b_1
X_3946_ _3946_/A vssd1 vssd1 vccd1 vccd1 _7542_/D sky130_fd_sc_hd__clkbuf_1
X_3877_ _3877_/A vssd1 vssd1 vccd1 vccd1 _7567_/D sky130_fd_sc_hd__clkbuf_1
X_5616_ _7091_/Q _5073_/A _5624_/S vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__mux2_1
X_6596_ _6534_/A _6604_/C _7511_/Q vssd1 vssd1 vccd1 vccd1 _6599_/B sky130_fd_sc_hd__a21o_1
X_5547_ _5547_/A vssd1 vssd1 vccd1 vccd1 _7065_/D sky130_fd_sc_hd__clkbuf_1
X_5478_ _5474_/X _7198_/Q input15/X _5475_/X vssd1 vssd1 vccd1 vccd1 _5478_/X sky130_fd_sc_hd__a22o_2
X_7217_ _7217_/CLK _7217_/D vssd1 vssd1 vccd1 vccd1 _7217_/Q sky130_fd_sc_hd__dfxtp_1
X_4429_ _4429_/A vssd1 vssd1 vccd1 vccd1 _7334_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3276_ _6670_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3276_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7148_ _7148_/CLK _7148_/D vssd1 vssd1 vccd1 vccd1 _7148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7079_ _7079_/CLK _7079_/D vssd1 vssd1 vccd1 vccd1 _7079_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__3111_ clkbuf_0__3111_/X vssd1 vssd1 vccd1 vccd1 _6437__68/A sky130_fd_sc_hd__clkbuf_16
XFILLER_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2757_ clkbuf_0__2757_/X vssd1 vssd1 vccd1 vccd1 _5810__299/A sky130_fd_sc_hd__clkbuf_16
XFILLER_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3800_ _3800_/A vssd1 vssd1 vccd1 vccd1 _7597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _7147_/Q _4340_/X _4782_/S vssd1 vssd1 vccd1 vccd1 _4781_/A sky130_fd_sc_hd__mux2_1
X_3731_ _4936_/A _3797_/C vssd1 vssd1 vccd1 vccd1 _3754_/S sky130_fd_sc_hd__nand2_2
XFILLER_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3662_ _3662_/A vssd1 vssd1 vccd1 vccd1 _7685_/D sky130_fd_sc_hd__clkbuf_1
X_6450_ _6450_/A _6450_/B vssd1 vssd1 vccd1 vccd1 _6451_/B sky130_fd_sc_hd__xnor2_1
X_3593_ _3593_/A vssd1 vssd1 vccd1 vccd1 _7703_/D sky130_fd_sc_hd__clkbuf_1
X_5401_ _5362_/S _7120_/Q _5252_/A vssd1 vssd1 vccd1 vccd1 _5401_/X sky130_fd_sc_hd__o21ba_1
X_5332_ _7546_/Q _5225_/X _5293_/A vssd1 vssd1 vccd1 vccd1 _5332_/X sky130_fd_sc_hd__o21ba_1
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5263_ _5363_/A _5259_/Y _5261_/Y _5396_/A vssd1 vssd1 vccd1 vccd1 _5263_/X sky130_fd_sc_hd__o211a_1
XFILLER_87_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4214_ _4236_/S vssd1 vssd1 vccd1 vccd1 _4227_/S sky130_fd_sc_hd__clkbuf_2
X_7002_ _7002_/A vssd1 vssd1 vccd1 vccd1 _7722_/D sky130_fd_sc_hd__clkbuf_1
X_5194_ _5481_/A _7061_/Q _5482_/A input3/X vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__a22o_1
X_4145_ _7437_/Q _3588_/X _4149_/S vssd1 vssd1 vccd1 vccd1 _4146_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4076_ _4175_/A _4642_/B vssd1 vssd1 vccd1 vccd1 _4092_/S sky130_fd_sc_hd__nor2_2
XFILLER_83_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4978_ _4978_/A vssd1 vssd1 vccd1 vccd1 _4978_/X sky130_fd_sc_hd__clkbuf_1
X_7697_ _7697_/CLK _7697_/D vssd1 vssd1 vccd1 vccd1 _7697_/Q sky130_fd_sc_hd__dfxtp_1
X_3929_ _4265_/B _4802_/A vssd1 vssd1 vccd1 vccd1 _3945_/S sky130_fd_sc_hd__or2_4
XFILLER_109_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6579_ _7507_/Q _6579_/B _6579_/C vssd1 vssd1 vccd1 vccd1 _6579_/Y sky130_fd_sc_hd__nand3_1
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6646__95 _6647__96/A vssd1 vssd1 vccd1 vccd1 _7539_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__2954_ clkbuf_0__2954_/X vssd1 vssd1 vccd1 vccd1 _6027__311/A sky130_fd_sc_hd__clkbuf_16
XFILLER_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _5901_/S _5943_/Y _5945_/Y _5947_/Y _5949_/Y vssd1 vssd1 vccd1 vccd1 _5950_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4901_ _4916_/S vssd1 vssd1 vccd1 vccd1 _4910_/S sky130_fd_sc_hd__buf_2
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7620_ _7620_/CLK _7620_/D vssd1 vssd1 vccd1 vccd1 _7620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5881_ _7219_/Q _5814_/X _5879_/X _5880_/X vssd1 vssd1 vccd1 vccd1 _7219_/D sky130_fd_sc_hd__o211a_1
XFILLER_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4832_ _4831_/X _7126_/Q _4835_/S vssd1 vssd1 vccd1 vccd1 _4833_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7551_ _7551_/CLK _7551_/D vssd1 vssd1 vccd1 vccd1 _7551_/Q sky130_fd_sc_hd__dfxtp_1
X_6653__101 _6656__104/A vssd1 vssd1 vccd1 vccd1 _7545_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__2630_ _5506_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2630_/X sky130_fd_sc_hd__clkbuf_16
X_4763_ _4763_/A vssd1 vssd1 vccd1 vccd1 _7156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7482_ _7482_/CLK _7482_/D vssd1 vssd1 vccd1 vccd1 _7482_/Q sky130_fd_sc_hd__dfxtp_1
X_3714_ _3469_/X _7629_/Q _3722_/S vssd1 vssd1 vccd1 vccd1 _3715_/A sky130_fd_sc_hd__mux2_1
X_4694_ _3819_/X _7210_/Q _4694_/S vssd1 vssd1 vccd1 vccd1 _4695_/A sky130_fd_sc_hd__mux2_1
X_6502_ _6469_/X _6470_/Y _6454_/A _6501_/Y _6454_/B vssd1 vssd1 vccd1 vccd1 _6504_/B
+ sky130_fd_sc_hd__a2111o_1
X_6433_ _6619_/A vssd1 vssd1 vccd1 vccd1 _6433_/X sky130_fd_sc_hd__buf_1
X_3645_ _3644_/X _7689_/Q _3657_/S vssd1 vssd1 vccd1 vccd1 _3646_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6364_ _6370_/A vssd1 vssd1 vccd1 vccd1 _6364_/X sky130_fd_sc_hd__buf_1
X_3576_ _4363_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _4364_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6295_ _6388_/A vssd1 vssd1 vccd1 vccd1 _6295_/X sky130_fd_sc_hd__buf_1
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5315_ _5315_/A _5315_/B vssd1 vssd1 vccd1 vccd1 _5315_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5246_ _7544_/Q _7434_/Q _7402_/Q _7386_/Q _5299_/A _4374_/A vssd1 vssd1 vccd1 vccd1
+ _5246_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5177_ _5360_/A _5174_/X _5176_/X _5163_/A vssd1 vssd1 vccd1 vccd1 _5177_/X sky130_fd_sc_hd__a211o_1
X_4128_ _4128_/A vssd1 vssd1 vccd1 vccd1 _7445_/D sky130_fd_sc_hd__clkbuf_1
X_4059_ _4074_/S vssd1 vssd1 vccd1 vccd1 _4068_/S sky130_fd_sc_hd__buf_2
X_6265__412 _6267__414/A vssd1 vssd1 vccd1 vccd1 _7352_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6717__153 _6718__154/A vssd1 vssd1 vccd1 vccd1 _7597_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3084_ clkbuf_0__3084_/X vssd1 vssd1 vccd1 vccd1 _6298__436/A sky130_fd_sc_hd__clkbuf_16
X_5100_ _5100_/A vssd1 vssd1 vccd1 vccd1 _5100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6080_ _6086_/A vssd1 vssd1 vccd1 vccd1 _6080_/X sky130_fd_sc_hd__buf_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A _5035_/B vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__and2_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6982_ _7275_/Q _7010_/B vssd1 vssd1 vccd1 vccd1 _7007_/S sky130_fd_sc_hd__nand2_2
X_5933_ _5882_/X _5918_/X _5932_/Y vssd1 vssd1 vccd1 vccd1 _5933_/X sky130_fd_sc_hd__a21o_1
X_5864_ _5862_/X _5863_/X _5959_/S vssd1 vssd1 vccd1 vccd1 _5864_/X sky130_fd_sc_hd__mux2_1
X_7603_ _7603_/CLK _7603_/D vssd1 vssd1 vccd1 vccd1 _7603_/Q sky130_fd_sc_hd__dfxtp_1
X_4815_ _4815_/A vssd1 vssd1 vccd1 vccd1 _7132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7534_ _7534_/CLK _7534_/D vssd1 vssd1 vccd1 vccd1 _7534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5795_ _5795_/A vssd1 vssd1 vccd1 vccd1 _7206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4746_ _7163_/Q _4340_/X _4748_/S vssd1 vssd1 vccd1 vccd1 _4747_/A sky130_fd_sc_hd__mux2_1
X_4677_ _4677_/A vssd1 vssd1 vccd1 vccd1 _7226_/D sky130_fd_sc_hd__clkbuf_1
X_7465_ _7465_/CLK _7465_/D vssd1 vssd1 vccd1 vccd1 _7465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7396_ _7396_/CLK _7396_/D vssd1 vssd1 vccd1 vccd1 _7396_/Q sky130_fd_sc_hd__dfxtp_1
X_3628_ _3542_/X _7692_/Q _3630_/S vssd1 vssd1 vccd1 vccd1 _3629_/A sky130_fd_sc_hd__mux2_1
X_6039__321 _6042__324/A vssd1 vssd1 vccd1 vccd1 _7247_/CLK sky130_fd_sc_hd__inv_2
X_3559_ _7347_/Q vssd1 vssd1 vccd1 vccd1 _4396_/A sky130_fd_sc_hd__inv_2
XFILLER_103_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5229_ _5381_/A _6274_/B vssd1 vssd1 vccd1 vccd1 _5308_/A sky130_fd_sc_hd__or2_2
XFILLER_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__3290_ clkbuf_0__3290_/X vssd1 vssd1 vccd1 vccd1 _6749__179/A sky130_fd_sc_hd__clkbuf_16
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2722_ clkbuf_0__2722_/X vssd1 vssd1 vccd1 vccd1 _5735__283/A sky130_fd_sc_hd__clkbuf_16
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4600_ _4255_/X _7260_/Q _4604_/S vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5580_ _5663_/A vssd1 vssd1 vccd1 vccd1 _5580_/X sky130_fd_sc_hd__buf_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4531_ _4531_/A vssd1 vssd1 vccd1 vccd1 _7291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7250_ _7250_/CLK _7250_/D vssd1 vssd1 vccd1 vccd1 _7250_/Q sky130_fd_sc_hd__dfxtp_1
X_4462_ _4462_/A vssd1 vssd1 vccd1 vccd1 _4477_/A sky130_fd_sc_hd__buf_4
X_6201_ _6201_/A vssd1 vssd1 vccd1 vccd1 _6201_/X sky130_fd_sc_hd__buf_1
XFILLER_98_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7181_ _7181_/CLK _7181_/D vssd1 vssd1 vccd1 vccd1 _7181_/Q sky130_fd_sc_hd__dfxtp_1
X_4393_ _5331_/A _4393_/B vssd1 vssd1 vccd1 vccd1 _4394_/C sky130_fd_sc_hd__nor2_1
X_6132_ _6121_/Y _6122_/X _6126_/Y _6130_/Y _6131_/X vssd1 vssd1 vccd1 vccd1 _6165_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5014_/A vssd1 vssd1 vccd1 vccd1 _5059_/A sky130_fd_sc_hd__buf_2
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5916_ _5914_/X _5915_/X _5998_/S vssd1 vssd1 vccd1 vccd1 _5916_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6342__472 _6342__472/A vssd1 vssd1 vccd1 vccd1 _7414_/CLK sky130_fd_sc_hd__inv_2
X_6896_ _7662_/Q _6892_/X _6895_/X _6880_/X vssd1 vssd1 vccd1 vccd1 _7661_/D sky130_fd_sc_hd__o211a_1
X_5847_ _4976_/A _3513_/X _6993_/A vssd1 vssd1 vccd1 vccd1 _6607_/A sky130_fd_sc_hd__a21o_4
XFILLER_22_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6969__1 _5499_/A vssd1 vssd1 vccd1 vccd1 _7711_/CLK sky130_fd_sc_hd__inv_2
X_5778_ _5022_/A _7199_/Q _5782_/S vssd1 vssd1 vccd1 vccd1 _5779_/A sky130_fd_sc_hd__mux2_1
X_7517_ _7517_/CLK _7517_/D vssd1 vssd1 vccd1 vccd1 _7517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4729_ _4729_/A vssd1 vssd1 vccd1 vccd1 _7171_/D sky130_fd_sc_hd__clkbuf_1
X_7448_ _7448_/CLK _7448_/D vssd1 vssd1 vccd1 vccd1 _7448_/Q sky130_fd_sc_hd__dfxtp_1
X_7379_ _7379_/CLK _7379_/D vssd1 vssd1 vccd1 vccd1 _7379_/Q sky130_fd_sc_hd__dfxtp_1
X_6666__111 _6666__111/A vssd1 vssd1 vccd1 vccd1 _7555_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6384__506 _6385__507/A vssd1 vssd1 vccd1 vccd1 _7448_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3273_ clkbuf_0__3273_/X vssd1 vssd1 vccd1 vccd1 _6664_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_25_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6020__306 _6021__307/A vssd1 vssd1 vccd1 vccd1 _7232_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5662__224 _5662__224/A vssd1 vssd1 vccd1 vccd1 _7118_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6285__426 _6288__429/A vssd1 vssd1 vccd1 vccd1 _7368_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6750_ _6938_/A vssd1 vssd1 vccd1 vccd1 _6750_/X sky130_fd_sc_hd__buf_1
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3962_ _3962_/A vssd1 vssd1 vccd1 vccd1 _7535_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__2636_ clkbuf_0__2636_/X vssd1 vssd1 vccd1 vccd1 _5523__194/A sky130_fd_sc_hd__clkbuf_16
X_3893_ _7560_/Q _3597_/X _3897_/S vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__mux2_1
X_5632_ _5632_/A vssd1 vssd1 vccd1 vccd1 _7098_/D sky130_fd_sc_hd__clkbuf_1
X_5563_ _7496_/Q vssd1 vssd1 vccd1 vccd1 _6610_/B sky130_fd_sc_hd__inv_2
XFILLER_117_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4514_ _7298_/Q _4331_/X _4516_/S vssd1 vssd1 vccd1 vccd1 _4515_/A sky130_fd_sc_hd__mux2_1
X_7302_ _7302_/CLK _7302_/D vssd1 vssd1 vccd1 vccd1 _7302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5494_ _7105_/Q _5493_/X _5494_/S vssd1 vssd1 vccd1 vccd1 _5495_/A sky130_fd_sc_hd__mux2_2
X_7233_ _7233_/CLK _7233_/D vssd1 vssd1 vccd1 vccd1 _7233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3292_ _6751_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3292_/X sky130_fd_sc_hd__clkbuf_16
X_4445_ _4445_/A _4445_/B vssd1 vssd1 vccd1 vccd1 _7318_/D sky130_fd_sc_hd__nor2_1
X_7164_ _7164_/CLK _7164_/D vssd1 vssd1 vccd1 vccd1 _7164_/Q sky130_fd_sc_hd__dfxtp_1
X_4376_ _3568_/X _4376_/B _4376_/C _4376_/D vssd1 vssd1 vccd1 vccd1 _4377_/B sky130_fd_sc_hd__and4b_1
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _6158_/A _6112_/A _6158_/B vssd1 vssd1 vccd1 vccd1 _6771_/A sky130_fd_sc_hd__a21oi_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7723_/CLK _7095_/D vssd1 vssd1 vccd1 vccd1 _7095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6879_ _7656_/Q _6879_/B _6879_/C vssd1 vssd1 vccd1 vccd1 _6879_/Y sky130_fd_sc_hd__nand3_1
XFILLER_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6390__510 _6392__512/A vssd1 vssd1 vccd1 vccd1 _7452_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6349__478 _6350__479/A vssd1 vssd1 vccd1 vccd1 _7420_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _4229_/X _7402_/Q _4236_/S vssd1 vssd1 vccd1 vccd1 _4231_/A sky130_fd_sc_hd__mux2_1
X_6252__403 _6252__403/A vssd1 vssd1 vccd1 vccd1 _7343_/CLK sky130_fd_sc_hd__inv_2
X_4161_ _4100_/X _7430_/Q _4167_/S vssd1 vssd1 vccd1 vccd1 _4162_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5523__194 _5523__194/A vssd1 vssd1 vccd1 vccd1 _7051_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6428__60 _6429__61/A vssd1 vssd1 vccd1 vccd1 _7482_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4092_ _7456_/Q _3819_/X _4092_/S vssd1 vssd1 vccd1 vccd1 _4093_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6802_ _7639_/Q _7638_/Q _7640_/Q vssd1 vssd1 vccd1 vccd1 _6819_/D sky130_fd_sc_hd__a21boi_2
XFILLER_24_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4994_ _4994_/A vssd1 vssd1 vccd1 vccd1 _4994_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3945_ _3668_/X _7542_/Q _3945_/S vssd1 vssd1 vccd1 vccd1 _3946_/A sky130_fd_sc_hd__mux2_1
X_6664_ _6664_/A vssd1 vssd1 vccd1 vccd1 _6664_/X sky130_fd_sc_hd__buf_1
X_3876_ _3750_/X _7567_/Q _3878_/S vssd1 vssd1 vccd1 vccd1 _3877_/A sky130_fd_sc_hd__mux2_1
X_5615_ _5637_/A vssd1 vssd1 vccd1 vccd1 _5624_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6595_ _6593_/X _6594_/X _6569_/X vssd1 vssd1 vccd1 vccd1 _7510_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5546_ _6917_/A _7065_/Q _5546_/S vssd1 vssd1 vccd1 vccd1 _5547_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5477_ _5474_/X _7197_/Q input13/X _5475_/X vssd1 vssd1 vccd1 vccd1 _5477_/X sky130_fd_sc_hd__a22o_2
X_7216_ _7216_/CLK _7216_/D vssd1 vssd1 vccd1 vccd1 _7216_/Q sky130_fd_sc_hd__dfxtp_1
X_4428_ _4226_/X _7334_/Q _4428_/S vssd1 vssd1 vccd1 vccd1 _4429_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3275_ _6664_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3275_/X sky130_fd_sc_hd__clkbuf_16
X_6192__372 _6194__374/A vssd1 vssd1 vccd1 vccd1 _7302_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4359_ _4301_/C _4361_/B _4358_/X vssd1 vssd1 vccd1 vccd1 _7354_/D sky130_fd_sc_hd__a21oi_1
X_7147_ _7147_/CLK _7147_/D vssd1 vssd1 vccd1 vccd1 _7147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7078_ _7078_/CLK _7078_/D vssd1 vssd1 vccd1 vccd1 _7078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5732__280 _5736__284/A vssd1 vssd1 vccd1 vccd1 _7174_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__3110_ clkbuf_0__3110_/X vssd1 vssd1 vccd1 vccd1 _6432__64/A sky130_fd_sc_hd__clkbuf_16
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6711__148 _6712__149/A vssd1 vssd1 vccd1 vccd1 _7592_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _3899_/A vssd1 vssd1 vccd1 vccd1 _3730_/X sky130_fd_sc_hd__buf_2
X_6397__516 _6399__518/A vssd1 vssd1 vccd1 vccd1 _7458_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3661_ _3660_/X _7685_/Q _3669_/S vssd1 vssd1 vccd1 vccd1 _3662_/A sky130_fd_sc_hd__mux2_1
X_3592_ _7703_/Q _3591_/X _3595_/S vssd1 vssd1 vccd1 vccd1 _3593_/A sky130_fd_sc_hd__mux2_1
X_5400_ _5291_/A _5397_/X _5399_/X _5413_/A vssd1 vssd1 vccd1 vccd1 _5400_/X sky130_fd_sc_hd__a211o_1
X_5331_ _5331_/A _5331_/B vssd1 vssd1 vccd1 vccd1 _5331_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7001_ _6981_/X _7001_/B vssd1 vssd1 vccd1 vccd1 _7002_/A sky130_fd_sc_hd__and2b_1
X_5262_ _5262_/A vssd1 vssd1 vccd1 vccd1 _5396_/A sky130_fd_sc_hd__clkbuf_2
X_4213_ _4864_/A _4265_/B vssd1 vssd1 vccd1 vccd1 _4236_/S sky130_fd_sc_hd__or2_2
X_5193_ _5450_/A vssd1 vssd1 vccd1 vccd1 _5482_/A sky130_fd_sc_hd__buf_4
XFILLER_110_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6033__316 _6035__318/A vssd1 vssd1 vccd1 vccd1 _7242_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4144_ _4144_/A vssd1 vssd1 vccd1 vccd1 _7438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4075_ _4075_/A vssd1 vssd1 vccd1 vccd1 _7464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6967__53 _6967__53/A vssd1 vssd1 vccd1 vccd1 _7709_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4977_ _6911_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__and2_1
X_7696_ _7696_/CLK _7696_/D vssd1 vssd1 vccd1 vccd1 _7696_/Q sky130_fd_sc_hd__dfxtp_1
X_6298__436 _6298__436/A vssd1 vssd1 vccd1 vccd1 _7378_/CLK sky130_fd_sc_hd__inv_2
X_3928_ _4846_/B vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__clkbuf_4
X_3859_ _3859_/A vssd1 vssd1 vccd1 vccd1 _7574_/D sky130_fd_sc_hd__clkbuf_1
X_6259__409 _6259__409/A vssd1 vssd1 vccd1 vccd1 _7349_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6578_ _6586_/C _6578_/B _6593_/C vssd1 vssd1 vccd1 vccd1 _6578_/X sky130_fd_sc_hd__or3b_1
XFILLER_59_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6422__55 _6424__57/A vssd1 vssd1 vccd1 vccd1 _7477_/CLK sky130_fd_sc_hd__inv_2
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6199__378 _6199__378/A vssd1 vssd1 vccd1 vccd1 _7308_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2953_ clkbuf_0__2953_/X vssd1 vssd1 vccd1 vccd1 _6049_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_77_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6405__523 _6406__524/A vssd1 vssd1 vccd1 vccd1 _7465_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4900_ _4900_/A _4918_/B vssd1 vssd1 vccd1 vccd1 _4916_/S sky130_fd_sc_hd__or2_2
X_5880_ _6599_/A vssd1 vssd1 vccd1 vccd1 _5880_/X sky130_fd_sc_hd__clkbuf_2
X_4831_ _7325_/Q vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__buf_2
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7550_ _7550_/CLK _7550_/D vssd1 vssd1 vccd1 vccd1 _7550_/Q sky130_fd_sc_hd__dfxtp_1
X_4762_ _4578_/X _7156_/Q _4766_/S vssd1 vssd1 vccd1 vccd1 _4763_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7481_ _7481_/CLK _7481_/D vssd1 vssd1 vccd1 vccd1 _7481_/Q sky130_fd_sc_hd__dfxtp_1
X_3713_ _3728_/S vssd1 vssd1 vccd1 vccd1 _3722_/S sky130_fd_sc_hd__buf_2
X_4693_ _4693_/A vssd1 vssd1 vccd1 vccd1 _7211_/D sky130_fd_sc_hd__clkbuf_1
X_6501_ _6507_/B _6507_/C _7504_/Q vssd1 vssd1 vccd1 vccd1 _6501_/Y sky130_fd_sc_hd__a21oi_1
X_3644_ _4566_/A vssd1 vssd1 vccd1 vccd1 _3644_/X sky130_fd_sc_hd__clkbuf_2
X_3575_ _5230_/A _5230_/B _5230_/C _5230_/D _7358_/Q vssd1 vssd1 vccd1 vccd1 _4363_/B
+ sky130_fd_sc_hd__o41a_2
X_5314_ _7530_/Q _7110_/Q _7562_/Q _7126_/Q _5148_/X _4382_/C vssd1 vssd1 vccd1 vccd1
+ _5315_/B sky130_fd_sc_hd__mux4_1
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3112_ _6439_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3112_/X sky130_fd_sc_hd__clkbuf_16
X_5245_ _5245_/A vssd1 vssd1 vccd1 vccd1 _5299_/A sky130_fd_sc_hd__buf_2
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5176_ _4396_/A _7138_/Q _5175_/X vssd1 vssd1 vccd1 vccd1 _5176_/X sky130_fd_sc_hd__o21a_1
X_6660__106 _6663__109/A vssd1 vssd1 vccd1 vccd1 _7550_/CLK sky130_fd_sc_hd__inv_2
X_4127_ _4103_/X _7445_/Q _4131_/S vssd1 vssd1 vccd1 vccd1 _4128_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4058_ _4175_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _4074_/S sky130_fd_sc_hd__or2b_2
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6306__443 _6307__444/A vssd1 vssd1 vccd1 vccd1 _7385_/CLK sky130_fd_sc_hd__inv_2
X_7679_ _7679_/CLK _7679_/D vssd1 vssd1 vccd1 vccd1 _7679_/Q sky130_fd_sc_hd__dfxtp_1
X_6079__349 _6079__349/A vssd1 vssd1 vccd1 vccd1 _7278_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6961__48 _6961__48/A vssd1 vssd1 vccd1 vccd1 _7704_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3083_ clkbuf_0__3083_/X vssd1 vssd1 vccd1 vccd1 _6308_/A sky130_fd_sc_hd__clkbuf_16
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5030_/X sky130_fd_sc_hd__clkbuf_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6724__158 _6724__158/A vssd1 vssd1 vccd1 vccd1 _7602_/CLK sky130_fd_sc_hd__inv_2
X_6981_ _7034_/A vssd1 vssd1 vccd1 vccd1 _6981_/X sky130_fd_sc_hd__clkbuf_1
X_5932_ _5902_/A _5931_/X _5833_/X vssd1 vssd1 vccd1 vccd1 _5932_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5863_ _7211_/Q _7037_/Q _7259_/Q _7251_/Q _5841_/X _4462_/A vssd1 vssd1 vccd1 vccd1
+ _5863_/X sky130_fd_sc_hd__mux4_2
X_7602_ _7602_/CLK _7602_/D vssd1 vssd1 vccd1 vccd1 _7602_/Q sky130_fd_sc_hd__dfxtp_1
X_4814_ _4578_/X _7132_/Q _4818_/S vssd1 vssd1 vccd1 vccd1 _4815_/A sky130_fd_sc_hd__mux2_1
X_5794_ _7206_/Q _5038_/A _5794_/S vssd1 vssd1 vccd1 vccd1 _5795_/A sky130_fd_sc_hd__mux2_1
X_7533_ _7533_/CLK _7533_/D vssd1 vssd1 vccd1 vccd1 _7533_/Q sky130_fd_sc_hd__dfxtp_2
X_4745_ _4745_/A vssd1 vssd1 vccd1 vccd1 _7164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__3419_ clkbuf_0__3419_/X vssd1 vssd1 vccd1 vccd1 _6950__39/A sky130_fd_sc_hd__clkbuf_16
X_4676_ _3819_/X _7226_/Q _4676_/S vssd1 vssd1 vccd1 vccd1 _4677_/A sky130_fd_sc_hd__mux2_1
X_7464_ _7464_/CLK _7464_/D vssd1 vssd1 vccd1 vccd1 _7464_/Q sky130_fd_sc_hd__dfxtp_1
X_7395_ _7395_/CLK _7395_/D vssd1 vssd1 vccd1 vccd1 _7395_/Q sky130_fd_sc_hd__dfxtp_1
X_3627_ _3627_/A vssd1 vssd1 vccd1 vccd1 _7693_/D sky130_fd_sc_hd__clkbuf_1
X_3558_ _3570_/C vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3489_ _7310_/Q _3822_/C vssd1 vssd1 vccd1 vccd1 _4466_/C sky130_fd_sc_hd__or2b_1
X_6277_ _6277_/A vssd1 vssd1 vccd1 vccd1 _6277_/X sky130_fd_sc_hd__buf_1
XFILLER_102_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5228_ _5219_/Y _5221_/Y _5224_/Y _5227_/Y _5433_/A vssd1 vssd1 vccd1 vccd1 _5228_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5159_ _5319_/A _5156_/X _5158_/X vssd1 vssd1 vccd1 vccd1 _5159_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6753__6 _6754__7/A vssd1 vssd1 vccd1 vccd1 _7625_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__2721_ clkbuf_0__2721_/X vssd1 vssd1 vccd1 vccd1 _5728__277/A sky130_fd_sc_hd__clkbuf_16
XFILLER_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6934__26 _6934__26/A vssd1 vssd1 vccd1 vccd1 _7682_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4530_ _4220_/X _7291_/Q _4534_/S vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__mux2_1
X_4461_ _5924_/A vssd1 vssd1 vccd1 vccd1 _4462_/A sky130_fd_sc_hd__buf_6
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7180_ _7180_/CLK _7180_/D vssd1 vssd1 vccd1 vccd1 _7180_/Q sky130_fd_sc_hd__dfxtp_1
X_6131_ _6821_/A _6452_/A _6452_/B vssd1 vssd1 vccd1 vccd1 _6131_/X sky130_fd_sc_hd__and3_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4392_ _5315_/A _4394_/B _4391_/Y vssd1 vssd1 vccd1 vccd1 _7349_/D sky130_fd_sc_hd__o21a_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6062_ _6086_/A vssd1 vssd1 vccd1 vccd1 _6062_/X sky130_fd_sc_hd__buf_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5013_/A vssd1 vssd1 vccd1 vccd1 _5013_/X sky130_fd_sc_hd__clkbuf_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5915_ _7245_/Q _7229_/Q _7475_/Q _7467_/Q _5860_/X _5861_/X vssd1 vssd1 vccd1 vccd1
+ _5915_/X sky130_fd_sc_hd__mux4_2
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6895_ _7661_/Q _6905_/B vssd1 vssd1 vccd1 vccd1 _6895_/X sky130_fd_sc_hd__or2_1
XFILLER_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5846_ _5902_/A _5846_/B vssd1 vssd1 vccd1 vccd1 _5846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5777_ _5777_/A vssd1 vssd1 vccd1 vccd1 _7198_/D sky130_fd_sc_hd__clkbuf_1
X_7516_ _7516_/CLK _7516_/D vssd1 vssd1 vccd1 vccd1 _7516_/Q sky130_fd_sc_hd__dfxtp_1
X_4728_ _4581_/X _7171_/Q _4730_/S vssd1 vssd1 vccd1 vccd1 _4729_/A sky130_fd_sc_hd__mux2_1
X_4659_ _4659_/A vssd1 vssd1 vccd1 vccd1 _7234_/D sky130_fd_sc_hd__clkbuf_1
X_7447_ _7447_/CLK _7447_/D vssd1 vssd1 vccd1 vccd1 _7447_/Q sky130_fd_sc_hd__dfxtp_1
X_7378_ _7378_/CLK _7378_/D vssd1 vssd1 vccd1 vccd1 _7378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3272_ clkbuf_0__3272_/X vssd1 vssd1 vccd1 vccd1 _6655__103/A sky130_fd_sc_hd__clkbuf_16
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3961_ _3920_/X _7535_/Q _3963_/S vssd1 vssd1 vccd1 vccd1 _3962_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5700_ _5700_/A vssd1 vssd1 vccd1 vccd1 _5700_/X sky130_fd_sc_hd__buf_1
X_3892_ _3892_/A vssd1 vssd1 vccd1 vccd1 _7561_/D sky130_fd_sc_hd__clkbuf_1
X_5631_ _7098_/Q _7197_/Q _5635_/S vssd1 vssd1 vccd1 vccd1 _5632_/A sky130_fd_sc_hd__mux2_1
X_5562_ _6561_/A vssd1 vssd1 vccd1 vccd1 _6579_/B sky130_fd_sc_hd__clkbuf_2
X_4513_ _4513_/A vssd1 vssd1 vccd1 vccd1 _7299_/D sky130_fd_sc_hd__clkbuf_1
X_7301_ _7301_/CLK _7301_/D vssd1 vssd1 vccd1 vccd1 _7301_/Q sky130_fd_sc_hd__dfxtp_1
X_7232_ _7232_/CLK _7232_/D vssd1 vssd1 vccd1 vccd1 _7232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5493_ _7080_/Q _5492_/X _5493_/S vssd1 vssd1 vccd1 vccd1 _5493_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3291_ _6750_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3291_/X sky130_fd_sc_hd__clkbuf_16
X_4444_ _4587_/B _4447_/A _4438_/X vssd1 vssd1 vccd1 vccd1 _4445_/B sky130_fd_sc_hd__o21ai_1
X_7163_ _7163_/CLK _7163_/D vssd1 vssd1 vccd1 vccd1 _7163_/Q sky130_fd_sc_hd__dfxtp_1
X_4375_ _4375_/A vssd1 vssd1 vccd1 vccd1 _5331_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _7723_/CLK _7094_/D vssd1 vssd1 vccd1 vccd1 _7094_/Q sky130_fd_sc_hd__dfxtp_1
X_6114_ _7655_/Q vssd1 vssd1 vccd1 vccd1 _6158_/B sky130_fd_sc_hd__inv_2
XFILLER_112_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6971__3 _6972__4/A vssd1 vssd1 vccd1 vccd1 _7713_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6878_ _6878_/A _6878_/B _6889_/B _6878_/D vssd1 vssd1 vccd1 vccd1 _6879_/C sky130_fd_sc_hd__or4_1
X_5829_ _5869_/A _5829_/B vssd1 vssd1 vccd1 vccd1 _5829_/X sky130_fd_sc_hd__or2_1
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6291__431 _6292__432/A vssd1 vssd1 vccd1 vccd1 _7373_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ _4160_/A vssd1 vssd1 vccd1 vccd1 _7431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4091_ _4091_/A vssd1 vssd1 vccd1 vccd1 _7457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6801_ _6794_/A _6781_/X _6886_/A _6794_/X _6800_/X vssd1 vssd1 vccd1 vccd1 _7639_/D
+ sky130_fd_sc_hd__o2111a_1
X_4993_ _4993_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _4994_/A sky130_fd_sc_hd__and2_1
X_6732_ _6732_/A vssd1 vssd1 vccd1 vccd1 _6732_/X sky130_fd_sc_hd__buf_1
X_3944_ _3944_/A vssd1 vssd1 vccd1 vccd1 _7543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3875_ _3875_/A vssd1 vssd1 vccd1 vccd1 _7568_/D sky130_fd_sc_hd__clkbuf_1
X_6761__13 _6761__13/A vssd1 vssd1 vccd1 vccd1 _7632_/CLK sky130_fd_sc_hd__inv_2
X_5614_ _5614_/A vssd1 vssd1 vccd1 vccd1 _7090_/D sky130_fd_sc_hd__clkbuf_1
X_6300__438 _6301__439/A vssd1 vssd1 vccd1 vccd1 _7380_/CLK sky130_fd_sc_hd__inv_2
X_6594_ _6594_/A _6609_/A _6594_/C vssd1 vssd1 vccd1 vccd1 _6594_/X sky130_fd_sc_hd__and3_1
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5545_ _5545_/A vssd1 vssd1 vccd1 vccd1 _7064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5476_ _5474_/X _7196_/Q input12/X _5475_/X vssd1 vssd1 vccd1 vccd1 _5476_/X sky130_fd_sc_hd__a22o_2
X_7215_ _7215_/CLK _7215_/D vssd1 vssd1 vccd1 vccd1 _7215_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3274_ _6658_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3274_/X sky130_fd_sc_hd__clkbuf_16
X_4427_ _4427_/A vssd1 vssd1 vccd1 vccd1 _7335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7146_ _7146_/CLK _7146_/D vssd1 vssd1 vccd1 vccd1 _7146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _3574_/A _4350_/B _4385_/A vssd1 vssd1 vccd1 vccd1 _4358_/X sky130_fd_sc_hd__a21o_1
X_4289_ _4246_/X _7381_/Q _4293_/S vssd1 vssd1 vccd1 vccd1 _4290_/A sky130_fd_sc_hd__mux2_1
X_7077_ _7077_/CLK _7077_/D vssd1 vssd1 vccd1 vccd1 _7077_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6355__483 _6355__483/A vssd1 vssd1 vccd1 vccd1 _7425_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_80 _6919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6679__122 _6680__123/A vssd1 vssd1 vccd1 vccd1 _7566_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3660_ _4578_/A vssd1 vssd1 vccd1 vccd1 _3660_/X sky130_fd_sc_hd__buf_2
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3591_ _7325_/Q vssd1 vssd1 vccd1 vccd1 _3591_/X sky130_fd_sc_hd__buf_4
X_5709__261 _5711__263/A vssd1 vssd1 vccd1 vccd1 _7155_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5330_ _7404_/Q _7388_/Q _5330_/S vssd1 vssd1 vccd1 vccd1 _5331_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7732_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5261_ _5360_/A _5261_/B vssd1 vssd1 vccd1 vccd1 _5261_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7000_ _4997_/A _6129_/A _7000_/S vssd1 vssd1 vccd1 vccd1 _7001_/B sky130_fd_sc_hd__mux2_1
X_4212_ _4900_/A vssd1 vssd1 vccd1 vccd1 _4864_/A sky130_fd_sc_hd__clkbuf_4
X_5192_ _5458_/A vssd1 vssd1 vccd1 vccd1 _5481_/A sky130_fd_sc_hd__buf_4
X_4143_ _7438_/Q _3585_/X _4149_/S vssd1 vssd1 vccd1 vccd1 _4144_/A sky130_fd_sc_hd__mux2_1
X_4074_ _3923_/X _7464_/Q _4074_/S vssd1 vssd1 vccd1 vccd1 _4075_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4976_ _4976_/A vssd1 vssd1 vccd1 vccd1 _6911_/A sky130_fd_sc_hd__clkbuf_16
X_7695_ _7695_/CLK _7695_/D vssd1 vssd1 vccd1 vccd1 _7695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3927_ _3927_/A _4363_/A _3927_/C vssd1 vssd1 vccd1 vccd1 _4846_/B sky130_fd_sc_hd__or3_4
X_3858_ _3753_/X _7574_/Q _3858_/S vssd1 vssd1 vccd1 vccd1 _3859_/A sky130_fd_sc_hd__mux2_1
X_3789_ _3789_/A vssd1 vssd1 vccd1 vccd1 _7600_/D sky130_fd_sc_hd__clkbuf_1
X_6577_ _7507_/Q _6577_/B vssd1 vssd1 vccd1 vccd1 _6578_/B sky130_fd_sc_hd__nor2_1
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5459_ _5458_/X _7190_/Q _5450_/X input6/X vssd1 vssd1 vccd1 vccd1 _5459_/X sky130_fd_sc_hd__a22o_1
X_5803__293 _5803__293/A vssd1 vssd1 vccd1 vccd1 _7211_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7129_ _7129_/CLK _7129_/D vssd1 vssd1 vccd1 vccd1 _7129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2952_ clkbuf_0__2952_/X vssd1 vssd1 vccd1 vccd1 _6021__307/A sky130_fd_sc_hd__clkbuf_16
XFILLER_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4830_ _4830_/A vssd1 vssd1 vccd1 vccd1 _7127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _4761_/A vssd1 vssd1 vccd1 vccd1 _7157_/D sky130_fd_sc_hd__clkbuf_1
X_7480_ _7480_/CLK _7480_/D vssd1 vssd1 vccd1 vccd1 _7480_/Q sky130_fd_sc_hd__dfxtp_1
X_3712_ _3797_/C _4678_/A vssd1 vssd1 vccd1 vccd1 _3728_/S sky130_fd_sc_hd__nand2_2
X_4692_ _3816_/X _7211_/Q _4694_/S vssd1 vssd1 vccd1 vccd1 _4693_/A sky130_fd_sc_hd__mux2_1
X_6500_ _6500_/A _6500_/B vssd1 vssd1 vccd1 vccd1 _6504_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3643_ _7327_/Q vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__clkbuf_4
X_5313_ _5481_/A _7065_/Q _5482_/A input29/X vssd1 vssd1 vccd1 vccd1 _5343_/A sky130_fd_sc_hd__a22oi_1
X_3574_ _3574_/A _4376_/D vssd1 vssd1 vccd1 vccd1 _5230_/D sky130_fd_sc_hd__and2_1
XFILLER_114_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3111_ _6433_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3111_/X sky130_fd_sc_hd__clkbuf_16
X_5244_ _7132_/Q _7055_/Q _7047_/Q _7268_/Q _5267_/A _5138_/X vssd1 vssd1 vccd1 vccd1
+ _5244_/X sky130_fd_sc_hd__mux4_1
X_5175_ _7517_/Q _5403_/S _5303_/A vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__o21ba_1
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _4126_/A vssd1 vssd1 vccd1 vccd1 _7446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4057_ _4057_/A vssd1 vssd1 vccd1 vccd1 _7472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ _5092_/A vssd1 vssd1 vccd1 vccd1 _4966_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__2757_ _5805_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2757_/X sky130_fd_sc_hd__clkbuf_16
X_7678_ _7678_/CLK _7678_/D vssd1 vssd1 vccd1 vccd1 _7678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6629_ _7525_/Q _6607_/A _6615_/A vssd1 vssd1 vccd1 vccd1 _7525_/D sky130_fd_sc_hd__a21o_1
XFILLER_106_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6946__35 _6948__37/A vssd1 vssd1 vccd1 vccd1 _7691_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3082_ clkbuf_0__3082_/X vssd1 vssd1 vccd1 vccd1 _6292__432/A sky130_fd_sc_hd__clkbuf_16
XFILLER_111_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6980_ _6980_/A vssd1 vssd1 vccd1 vccd1 _7716_/D sky130_fd_sc_hd__clkbuf_1
X_5931_ _5901_/S _5920_/Y _5923_/Y _5927_/Y _5930_/Y vssd1 vssd1 vccd1 vccd1 _5931_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6368__493 _6368__493/A vssd1 vssd1 vccd1 vccd1 _7435_/CLK sky130_fd_sc_hd__inv_2
X_5862_ _7243_/Q _7227_/Q _7473_/Q _7465_/Q _5860_/X _5861_/X vssd1 vssd1 vccd1 vccd1
+ _5862_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7601_ _7601_/CLK _7601_/D vssd1 vssd1 vccd1 vccd1 _7601_/Q sky130_fd_sc_hd__dfxtp_1
X_4813_ _4813_/A vssd1 vssd1 vccd1 vccd1 _7133_/D sky130_fd_sc_hd__clkbuf_1
X_5793_ _5793_/A vssd1 vssd1 vccd1 vccd1 _7205_/D sky130_fd_sc_hd__clkbuf_1
X_7532_ _7532_/CLK _7532_/D vssd1 vssd1 vccd1 vccd1 _7532_/Q sky130_fd_sc_hd__dfxtp_2
X_4744_ _7164_/Q _4337_/X _4748_/S vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__3418_ clkbuf_0__3418_/X vssd1 vssd1 vccd1 vccd1 _6941__31/A sky130_fd_sc_hd__clkbuf_16
X_4675_ _4675_/A vssd1 vssd1 vccd1 vccd1 _7227_/D sky130_fd_sc_hd__clkbuf_1
X_7463_ _7463_/CLK _7463_/D vssd1 vssd1 vccd1 vccd1 _7463_/Q sky130_fd_sc_hd__dfxtp_1
X_7394_ _7394_/CLK _7394_/D vssd1 vssd1 vccd1 vccd1 _7394_/Q sky130_fd_sc_hd__dfxtp_1
X_3626_ _3538_/X _7693_/Q _3630_/S vssd1 vssd1 vccd1 vccd1 _3627_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6345_ _6351_/A vssd1 vssd1 vccd1 vccd1 _6345_/X sky130_fd_sc_hd__buf_1
X_3557_ _7352_/Q vssd1 vssd1 vccd1 vccd1 _3570_/C sky130_fd_sc_hd__clkbuf_1
X_3488_ _7318_/Q _3485_/Y _4443_/A _4467_/B vssd1 vssd1 vccd1 vccd1 _3493_/A sky130_fd_sc_hd__o211a_1
X_5227_ _5257_/A _5226_/X _5205_/X vssd1 vssd1 vccd1 vccd1 _5227_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_102_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5158_ _5178_/A vssd1 vssd1 vccd1 vccd1 _5158_/X sky130_fd_sc_hd__clkbuf_2
X_5089_ _5089_/A vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4109_ _7670_/Q vssd1 vssd1 vccd1 vccd1 _4109_/X sky130_fd_sc_hd__buf_2
XFILLER_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6046__327 _6046__327/A vssd1 vssd1 vccd1 vccd1 _7253_/CLK sky130_fd_sc_hd__inv_2
X_6085__354 _6085__354/A vssd1 vssd1 vccd1 vccd1 _7283_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2720_ clkbuf_0__2720_/X vssd1 vssd1 vccd1 vccd1 _5723__273/A sky130_fd_sc_hd__clkbuf_16
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _7311_/Q vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__clkbuf_2
X_6730__163 _6731__164/A vssd1 vssd1 vccd1 vccd1 _7607_/CLK sky130_fd_sc_hd__inv_2
X_4391_ _6274_/A _4391_/B vssd1 vssd1 vccd1 vccd1 _4391_/Y sky130_fd_sc_hd__nor2_1
X_6130_ _6777_/A _6789_/A vssd1 vssd1 vccd1 vccd1 _6130_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5012_/A _5012_/B vssd1 vssd1 vccd1 vccd1 _5013_/A sky130_fd_sc_hd__and2_1
XFILLER_112_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6963_ _6963_/A vssd1 vssd1 vccd1 vccd1 _6963_/X sky130_fd_sc_hd__buf_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5914_ _7213_/Q _7039_/Q _7261_/Q _7253_/Q _5912_/X _5913_/X vssd1 vssd1 vccd1 vccd1
+ _5914_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6894_ _7661_/Q _6892_/X _6893_/X _6880_/X vssd1 vssd1 vccd1 vccd1 _7660_/D sky130_fd_sc_hd__o211a_1
X_5845_ _5840_/X _5844_/X _5917_/A vssd1 vssd1 vccd1 vccd1 _5846_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5776_ _5020_/A _7198_/Q _5776_/S vssd1 vssd1 vccd1 vccd1 _5777_/A sky130_fd_sc_hd__mux2_1
X_7515_ _7516_/CLK _7515_/D vssd1 vssd1 vccd1 vccd1 _7515_/Q sky130_fd_sc_hd__dfxtp_1
X_4727_ _4727_/A vssd1 vssd1 vccd1 vccd1 _7172_/D sky130_fd_sc_hd__clkbuf_1
X_6418__534 _6418__534/A vssd1 vssd1 vccd1 vccd1 _7476_/CLK sky130_fd_sc_hd__inv_2
X_4658_ _4261_/X _7234_/Q _4658_/S vssd1 vssd1 vccd1 vccd1 _4659_/A sky130_fd_sc_hd__mux2_1
X_7446_ _7446_/CLK _7446_/D vssd1 vssd1 vccd1 vccd1 _7446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3609_ _3609_/A vssd1 vssd1 vccd1 vccd1 _3796_/C sky130_fd_sc_hd__clkbuf_2
Xinput90 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _5555_/A sky130_fd_sc_hd__buf_4
X_4589_ _4604_/S vssd1 vssd1 vccd1 vccd1 _4598_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7377_ _7377_/CLK _7377_/D vssd1 vssd1 vccd1 vccd1 _7377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3271_ clkbuf_0__3271_/X vssd1 vssd1 vccd1 vccd1 _6647__96/A sky130_fd_sc_hd__clkbuf_16
X_6673__117 _6675__119/A vssd1 vssd1 vccd1 vccd1 _7561_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6319__454 _6319__454/A vssd1 vssd1 vccd1 vccd1 _7396_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3960_ _3960_/A vssd1 vssd1 vccd1 vccd1 _7536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3891_ _7561_/Q _3594_/X _3891_/S vssd1 vssd1 vccd1 vccd1 _3892_/A sky130_fd_sc_hd__mux2_1
X_5630_ _5630_/A vssd1 vssd1 vccd1 vccd1 _7097_/D sky130_fd_sc_hd__clkbuf_1
X_5561_ _7497_/Q vssd1 vssd1 vccd1 vccd1 _6561_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5492_ _5492_/A input2/X vssd1 vssd1 vccd1 vccd1 _5492_/X sky130_fd_sc_hd__or2_4
XFILLER_117_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4512_ _7299_/Q _4328_/X _4516_/S vssd1 vssd1 vccd1 vccd1 _4513_/A sky130_fd_sc_hd__mux2_1
X_7300_ _7300_/CLK _7300_/D vssd1 vssd1 vccd1 vccd1 _7300_/Q sky130_fd_sc_hd__dfxtp_1
X_7231_ _7231_/CLK _7231_/D vssd1 vssd1 vccd1 vccd1 _7231_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3290_ _6744_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3290_/X sky130_fd_sc_hd__clkbuf_16
X_4443_ _4443_/A _4443_/B vssd1 vssd1 vccd1 vccd1 _4447_/A sky130_fd_sc_hd__and2_1
X_4374_ _4374_/A vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__buf_2
X_7162_ _7162_/CLK _7162_/D vssd1 vssd1 vccd1 vccd1 _7162_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7723_/CLK _7093_/D vssd1 vssd1 vccd1 vccd1 _7093_/Q sky130_fd_sc_hd__dfxtp_1
X_6113_ _6463_/A vssd1 vssd1 vccd1 vccd1 _6158_/A sky130_fd_sc_hd__inv_2
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6877_ _6794_/A _6878_/D _6781_/A vssd1 vssd1 vccd1 vccd1 _6879_/B sky130_fd_sc_hd__a21oi_2
X_6737__169 _6737__169/A vssd1 vssd1 vccd1 vccd1 _7613_/CLK sky130_fd_sc_hd__inv_2
X_5828_ _7408_/Q _7376_/Q _7707_/Q _7630_/Q _5921_/A _5856_/A vssd1 vssd1 vccd1 vccd1
+ _5829_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5759_ _5759_/A vssd1 vssd1 vccd1 vccd1 _7190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7429_ _7429_/CLK _7429_/D vssd1 vssd1 vccd1 vccd1 _7429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6059__337 _6060__338/A vssd1 vssd1 vccd1 vccd1 _7263_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4090_ _7457_/Q _3816_/X _4092_/S vssd1 vssd1 vccd1 vccd1 _4091_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ _6800_/A _6803_/B _6781_/X vssd1 vssd1 vccd1 vccd1 _6800_/X sky130_fd_sc_hd__or3b_1
X_4992_ _5106_/B vssd1 vssd1 vccd1 vccd1 _5001_/B sky130_fd_sc_hd__clkbuf_1
X_3943_ _3664_/X _7543_/Q _3945_/S vssd1 vssd1 vccd1 vccd1 _3944_/A sky130_fd_sc_hd__mux2_1
X_3874_ _3747_/X _7568_/Q _3878_/S vssd1 vssd1 vccd1 vccd1 _3875_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5613_ _7090_/Q _5071_/A _5613_/S vssd1 vssd1 vccd1 vccd1 _5614_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6593_ _6604_/C _6593_/B _6593_/C vssd1 vssd1 vccd1 vccd1 _6593_/X sky130_fd_sc_hd__and3b_1
X_5544_ _6915_/A _7064_/Q _5546_/S vssd1 vssd1 vccd1 vccd1 _5545_/A sky130_fd_sc_hd__mux2_1
X_5475_ _5482_/A vssd1 vssd1 vccd1 vccd1 _5475_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7214_ _7214_/CLK _7214_/D vssd1 vssd1 vccd1 vccd1 _7214_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3273_ _6657_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3273_/X sky130_fd_sc_hd__clkbuf_16
X_4426_ _4223_/X _7335_/Q _4428_/S vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__mux2_1
X_7145_ _7145_/CLK _7145_/D vssd1 vssd1 vccd1 vccd1 _7145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _4357_/A vssd1 vssd1 vccd1 vccd1 _7355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4288_ _4288_/A vssd1 vssd1 vccd1 vccd1 _7382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7076_ _7076_/CLK _7076_/D vssd1 vssd1 vccd1 vccd1 _7076_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6434__65 _6437__68/A vssd1 vssd1 vccd1 vccd1 _7487_/CLK sky130_fd_sc_hd__inv_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_70 _7306_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_81 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6362__488 _6363__489/A vssd1 vssd1 vccd1 vccd1 _7430_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3590_ _3590_/A vssd1 vssd1 vccd1 vccd1 _7704_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__3099_ clkbuf_0__3099_/X vssd1 vssd1 vccd1 vccd1 _6381__504/A sky130_fd_sc_hd__clkbuf_16
X_5260_ _7685_/Q _7608_/Q _5391_/S vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4211_ _4560_/A vssd1 vssd1 vccd1 vccd1 _4211_/X sky130_fd_sc_hd__buf_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5191_ _5191_/A vssd1 vssd1 vccd1 vccd1 _5458_/A sky130_fd_sc_hd__clkbuf_2
X_4142_ _4142_/A vssd1 vssd1 vccd1 vccd1 _7439_/D sky130_fd_sc_hd__clkbuf_1
X_4073_ _4073_/A vssd1 vssd1 vccd1 vccd1 _7465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4975_ _4975_/A vssd1 vssd1 vccd1 vccd1 _4975_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3926_ _3926_/A _4301_/C _3983_/B vssd1 vssd1 vccd1 vccd1 _4265_/B sky130_fd_sc_hd__or3b_4
X_7694_ _7694_/CLK _7694_/D vssd1 vssd1 vccd1 vccd1 _7694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3857_ _3857_/A vssd1 vssd1 vccd1 vccd1 _7575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6645_ _6645_/A vssd1 vssd1 vccd1 vccd1 _6645_/X sky130_fd_sc_hd__buf_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3788_ _3747_/X _7600_/Q _3792_/S vssd1 vssd1 vccd1 vccd1 _3789_/A sky130_fd_sc_hd__mux2_1
X_6576_ _7507_/Q _7506_/Q _7505_/Q _6576_/D vssd1 vssd1 vccd1 vccd1 _6586_/C sky130_fd_sc_hd__and4_1
XFILLER_118_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_193 vssd1 vssd1 vccd1 vccd1 CaravelHost_193/HI core0Index[0] sky130_fd_sc_hd__conb_1
X_5458_ _5458_/A vssd1 vssd1 vccd1 vccd1 _5458_/X sky130_fd_sc_hd__clkbuf_2
X_5389_ _7548_/Q _5290_/S _5303_/X vssd1 vssd1 vccd1 vccd1 _5389_/X sky130_fd_sc_hd__o21ba_1
X_4409_ _4409_/A vssd1 vssd1 vccd1 vccd1 _7343_/D sky130_fd_sc_hd__clkbuf_1
X_7128_ _7128_/CLK _7128_/D vssd1 vssd1 vccd1 vccd1 _7128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7059_ _7059_/CLK _7059_/D vssd1 vssd1 vccd1 vccd1 _7059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2951_ clkbuf_0__2951_/X vssd1 vssd1 vccd1 vccd1 _6015__302/A sky130_fd_sc_hd__clkbuf_16
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4760_ _4575_/X _7157_/Q _4760_/S vssd1 vssd1 vccd1 vccd1 _4761_/A sky130_fd_sc_hd__mux2_1
X_4691_ _4691_/A vssd1 vssd1 vccd1 vccd1 _7212_/D sky130_fd_sc_hd__clkbuf_1
X_3711_ _3861_/C _4436_/A _3711_/C vssd1 vssd1 vccd1 vccd1 _4678_/A sky130_fd_sc_hd__and3b_4
X_3642_ _3642_/A vssd1 vssd1 vccd1 vccd1 _7690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5312_ _5312_/A vssd1 vssd1 vccd1 vccd1 _5312_/X sky130_fd_sc_hd__clkbuf_1
X_3573_ _3573_/A _3573_/B vssd1 vssd1 vccd1 vccd1 _5230_/C sky130_fd_sc_hd__nand2_1
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6412__529 _6412__529/A vssd1 vssd1 vccd1 vccd1 _7471_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3110_ _6427_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3110_/X sky130_fd_sc_hd__clkbuf_16
X_5243_ _7348_/Q vssd1 vssd1 vccd1 vccd1 _5267_/A sky130_fd_sc_hd__buf_2
XFILLER_102_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5174_ _7154_/Q _7146_/Q _5285_/S vssd1 vssd1 vccd1 vccd1 _5174_/X sky130_fd_sc_hd__mux2_1
X_4125_ _4100_/X _7446_/Q _4131_/S vssd1 vssd1 vccd1 vccd1 _4126_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4056_ _3923_/X _7472_/Q _4056_/S vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4958_ _5014_/A vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3909_ _3908_/X _7555_/Q _3915_/S vssd1 vssd1 vccd1 vccd1 _3910_/A sky130_fd_sc_hd__mux2_1
X_7677_ _7677_/CLK _7677_/D vssd1 vssd1 vccd1 vccd1 _7677_/Q sky130_fd_sc_hd__dfxtp_1
X_4889_ _4889_/A vssd1 vssd1 vccd1 vccd1 _7077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6559_ _6562_/A _6559_/B vssd1 vssd1 vccd1 vccd1 _6560_/B sky130_fd_sc_hd__or2_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6313__449 _6313__449/A vssd1 vssd1 vccd1 vccd1 _7391_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5658__220 _5662__224/A vssd1 vssd1 vccd1 vccd1 _7114_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3081_ clkbuf_0__3081_/X vssd1 vssd1 vccd1 vccd1 _6288__429/A sky130_fd_sc_hd__clkbuf_16
XFILLER_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5930_ _5888_/A _5928_/X _5929_/X vssd1 vssd1 vccd1 vccd1 _5930_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5861_ _5870_/A vssd1 vssd1 vccd1 vccd1 _5861_/X sky130_fd_sc_hd__buf_2
X_7600_ _7600_/CLK _7600_/D vssd1 vssd1 vccd1 vccd1 _7600_/Q sky130_fd_sc_hd__dfxtp_1
X_4812_ _4575_/X _7133_/Q _4812_/S vssd1 vssd1 vccd1 vccd1 _4813_/A sky130_fd_sc_hd__mux2_1
X_5792_ _7205_/Q _5035_/A _5794_/S vssd1 vssd1 vccd1 vccd1 _5793_/A sky130_fd_sc_hd__mux2_1
X_7531_ _7531_/CLK _7531_/D vssd1 vssd1 vccd1 vccd1 _7531_/Q sky130_fd_sc_hd__dfxtp_1
X_4743_ _4743_/A vssd1 vssd1 vccd1 vccd1 _7165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7462_ _7462_/CLK _7462_/D vssd1 vssd1 vccd1 vccd1 _7462_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__3417_ clkbuf_0__3417_/X vssd1 vssd1 vccd1 vccd1 _6951_/A sky130_fd_sc_hd__clkbuf_16
X_4674_ _3816_/X _7227_/Q _4676_/S vssd1 vssd1 vccd1 vccd1 _4675_/A sky130_fd_sc_hd__mux2_1
X_6413_ _6413_/A vssd1 vssd1 vccd1 vccd1 _6413_/X sky130_fd_sc_hd__buf_1
X_7393_ _7393_/CLK _7393_/D vssd1 vssd1 vccd1 vccd1 _7393_/Q sky130_fd_sc_hd__dfxtp_1
X_3625_ _3625_/A vssd1 vssd1 vccd1 vccd1 _7694_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__3279_ clkbuf_0__3279_/X vssd1 vssd1 vccd1 vccd1 _6701_/A sky130_fd_sc_hd__clkbuf_16
X_3556_ _7353_/Q vssd1 vssd1 vccd1 vccd1 _3927_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3487_ _7318_/Q _3485_/Y _4443_/A _4467_/B vssd1 vssd1 vccd1 vccd1 _3494_/C sky130_fd_sc_hd__a31o_1
X_5226_ _7131_/Q _7054_/Q _7046_/Q _7267_/Q _5207_/X _5225_/X vssd1 vssd1 vccd1 vccd1
+ _5226_/X sky130_fd_sc_hd__mux4_1
X_5503__183 _5504__184/A vssd1 vssd1 vccd1 vccd1 _7039_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5157_ _7350_/Q vssd1 vssd1 vccd1 vccd1 _5178_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5088_ _7197_/Q _5090_/B vssd1 vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__and2_1
X_4108_ _4108_/A vssd1 vssd1 vccd1 vccd1 _7452_/D sky130_fd_sc_hd__clkbuf_1
X_4039_ _4587_/C _4587_/B _4039_/C vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__and3_2
XFILLER_112_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7729_ _7731_/CLK _7729_/D vssd1 vssd1 vccd1 vccd1 _7729_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5519__190 _5522__193/A vssd1 vssd1 vccd1 vccd1 _7047_/CLK sky130_fd_sc_hd__inv_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4390_ _5331_/A _4393_/B vssd1 vssd1 vccd1 vccd1 _4394_/B sky130_fd_sc_hd__and2_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5011_/A vssd1 vssd1 vccd1 vccd1 _5011_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5913_ _5924_/A vssd1 vssd1 vccd1 vccd1 _5913_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6893_ _7660_/Q _6893_/B vssd1 vssd1 vccd1 vccd1 _6893_/X sky130_fd_sc_hd__or2_1
X_5844_ _5842_/X _5843_/X _5910_/A vssd1 vssd1 vccd1 vccd1 _5844_/X sky130_fd_sc_hd__mux2_1
X_6630__82 _6632__84/A vssd1 vssd1 vccd1 vccd1 _7526_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7514_ _7516_/CLK _7514_/D vssd1 vssd1 vccd1 vccd1 _7514_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5775_ _5775_/A vssd1 vssd1 vccd1 vccd1 _7197_/D sky130_fd_sc_hd__clkbuf_1
X_4726_ _4578_/X _7172_/Q _4730_/S vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__mux2_1
X_4657_ _4657_/A vssd1 vssd1 vccd1 vccd1 _7235_/D sky130_fd_sc_hd__clkbuf_1
X_7445_ _7445_/CLK _7445_/D vssd1 vssd1 vccd1 vccd1 _7445_/Q sky130_fd_sc_hd__dfxtp_1
X_3608_ _4095_/B _4039_/C _4587_/C vssd1 vssd1 vccd1 vccd1 _4542_/B sky130_fd_sc_hd__and3b_2
Xinput80 wbs_data_i[4] vssd1 vssd1 vccd1 vccd1 _6917_/A sky130_fd_sc_hd__buf_8
Xinput91 wbs_we_i vssd1 vssd1 vccd1 vccd1 _5642_/A sky130_fd_sc_hd__buf_6
X_7376_ _7376_/CLK _7376_/D vssd1 vssd1 vccd1 vccd1 _7376_/Q sky130_fd_sc_hd__dfxtp_1
X_4588_ _4660_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4604_/S sky130_fd_sc_hd__nand2_2
X_6327_ _6333_/A vssd1 vssd1 vccd1 vccd1 _6327_/X sky130_fd_sc_hd__buf_1
X_3539_ _3538_/X _7709_/Q _3547_/S vssd1 vssd1 vccd1 vccd1 _3540_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6052__332 _6052__332/A vssd1 vssd1 vccd1 vccd1 _7258_/CLK sky130_fd_sc_hd__inv_2
X_5209_ _4396_/X _7139_/Q _5208_/X vssd1 vssd1 vccd1 vccd1 _5209_/X sky130_fd_sc_hd__o21a_1
X_6189_ _6195_/A vssd1 vssd1 vccd1 vccd1 _6189_/X sky130_fd_sc_hd__buf_1
XFILLER_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3270_ clkbuf_0__3270_/X vssd1 vssd1 vccd1 vccd1 _6644__94/A sky130_fd_sc_hd__clkbuf_16
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6243__395 _6246__398/A vssd1 vssd1 vccd1 vccd1 _7335_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5703__257 _5705__259/A vssd1 vssd1 vccd1 vccd1 _7151_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3890_ _3890_/A vssd1 vssd1 vccd1 vccd1 _7562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _7070_/Q _7069_/Q _5645_/A _5557_/X vssd1 vssd1 vccd1 vccd1 _7070_/D sky130_fd_sc_hd__o31a_1
XFILLER_117_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4511_ _4511_/A vssd1 vssd1 vccd1 vccd1 _7300_/D sky130_fd_sc_hd__clkbuf_1
X_5491_ _5375_/X _7209_/Q input27/X _5376_/X vssd1 vssd1 vccd1 vccd1 _5491_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7230_ _7230_/CLK _7230_/D vssd1 vssd1 vccd1 vccd1 _7230_/Q sky130_fd_sc_hd__dfxtp_1
X_4442_ _4587_/C _4445_/A _4441_/Y vssd1 vssd1 vccd1 vccd1 _7319_/D sky130_fd_sc_hd__o21a_1
XFILLER_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4373_ _5303_/A vssd1 vssd1 vccd1 vccd1 _4374_/A sky130_fd_sc_hd__clkbuf_2
X_7161_ _7161_/CLK _7161_/D vssd1 vssd1 vccd1 vccd1 _7161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6112_/A _6792_/A vssd1 vssd1 vccd1 vccd1 _6778_/A sky130_fd_sc_hd__xnor2_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7723_/CLK _7092_/D vssd1 vssd1 vccd1 vccd1 _7092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6043_ _6049_/A vssd1 vssd1 vccd1 vccd1 _6043_/X sky130_fd_sc_hd__buf_1
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6945_ _6963_/A vssd1 vssd1 vccd1 vccd1 _6945_/X sky130_fd_sc_hd__buf_1
XFILLER_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6876_ _6876_/A vssd1 vssd1 vccd1 vccd1 _6893_/B sky130_fd_sc_hd__clkbuf_2
X_5827_ _7311_/Q vssd1 vssd1 vccd1 vccd1 _5921_/A sky130_fd_sc_hd__buf_2
X_5758_ _5001_/A _7190_/Q _5758_/S vssd1 vssd1 vccd1 vccd1 _5759_/A sky130_fd_sc_hd__mux2_1
X_4709_ _4709_/A vssd1 vssd1 vccd1 vccd1 _7180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7428_ _7428_/CLK _7428_/D vssd1 vssd1 vccd1 vccd1 _7428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7359_ _7359_/CLK _7359_/D vssd1 vssd1 vccd1 vccd1 _7359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4991_ _4991_/A vssd1 vssd1 vccd1 vccd1 _4991_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _3942_/A vssd1 vssd1 vccd1 vccd1 _7544_/D sky130_fd_sc_hd__clkbuf_1
X_3873_ _3873_/A vssd1 vssd1 vccd1 vccd1 _7569_/D sky130_fd_sc_hd__clkbuf_1
X_5612_ _5612_/A vssd1 vssd1 vccd1 vccd1 _7089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6592_ _6594_/A _6592_/B vssd1 vssd1 vccd1 vccd1 _6593_/B sky130_fd_sc_hd__or2_1
X_5543_ _5543_/A vssd1 vssd1 vccd1 vccd1 _7063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5474_ _5481_/A vssd1 vssd1 vccd1 vccd1 _5474_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7213_ _7213_/CLK _7213_/D vssd1 vssd1 vccd1 vccd1 _7213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3272_ _6651_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3272_/X sky130_fd_sc_hd__clkbuf_16
X_4425_ _4425_/A vssd1 vssd1 vccd1 vccd1 _7336_/D sky130_fd_sc_hd__clkbuf_1
X_4356_ _6272_/C _4356_/B _4356_/C vssd1 vssd1 vccd1 vccd1 _4357_/A sky130_fd_sc_hd__and3_1
X_7144_ _7144_/CLK _7144_/D vssd1 vssd1 vccd1 vccd1 _7144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4287_ _4243_/X _7382_/Q _4293_/S vssd1 vssd1 vccd1 vccd1 _4288_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7075_ _7075_/CLK _7075_/D vssd1 vssd1 vccd1 vccd1 _7075_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6743__174 _6743__174/A vssd1 vssd1 vccd1 vccd1 _7618_/CLK sky130_fd_sc_hd__inv_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5652__215 _5655__218/A vssd1 vssd1 vccd1 vccd1 _7109_/CLK sky130_fd_sc_hd__inv_2
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6859_ _6857_/X _6859_/B _6859_/C vssd1 vssd1 vccd1 vccd1 _6860_/A sky130_fd_sc_hd__and3b_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_60 _3920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_71 _7309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_82 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6065__342 _6065__342/A vssd1 vssd1 vccd1 vccd1 _7268_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__3098_ clkbuf_0__3098_/X vssd1 vssd1 vccd1 vccd1 _6375__499/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6686__128 _6687__129/A vssd1 vssd1 vccd1 vccd1 _7572_/CLK sky130_fd_sc_hd__inv_2
X_4210_ _4210_/A vssd1 vssd1 vccd1 vccd1 _7408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5190_ _7732_/Q _5469_/C _5129_/Y _5189_/X vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__a22o_1
X_4141_ _7439_/Q _3549_/X _4149_/S vssd1 vssd1 vccd1 vccd1 _4142_/A sky130_fd_sc_hd__mux2_1
X_4072_ _3920_/X _7465_/Q _4074_/S vssd1 vssd1 vccd1 vccd1 _4073_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5716__267 _5716__267/A vssd1 vssd1 vccd1 vccd1 _7161_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4974_ _6908_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4975_/A sky130_fd_sc_hd__and2_1
XFILLER_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6713_ _6713_/A vssd1 vssd1 vccd1 vccd1 _6713_/X sky130_fd_sc_hd__buf_1
X_3925_ _3925_/A vssd1 vssd1 vccd1 vccd1 _7550_/D sky130_fd_sc_hd__clkbuf_1
X_7693_ _7693_/CLK _7693_/D vssd1 vssd1 vccd1 vccd1 _7693_/Q sky130_fd_sc_hd__dfxtp_1
X_3856_ _3750_/X _7575_/Q _3858_/S vssd1 vssd1 vccd1 vccd1 _3857_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3787_ _3787_/A vssd1 vssd1 vccd1 vccd1 _7601_/D sky130_fd_sc_hd__clkbuf_1
X_6575_ _6573_/Y _6574_/X _6569_/X vssd1 vssd1 vccd1 vccd1 _7506_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5457_ _7721_/Q _5448_/X _5449_/X _5456_/X vssd1 vssd1 vccd1 vccd1 _5457_/X sky130_fd_sc_hd__a31o_1
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XCaravelHost_194 vssd1 vssd1 vccd1 vccd1 CaravelHost_194/HI core0Index[1] sky130_fd_sc_hd__conb_1
X_4408_ _7343_/Q _4331_/X _4410_/S vssd1 vssd1 vccd1 vccd1 _4409_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5388_ _7136_/Q _7059_/Q _7051_/Q _7272_/Q _4374_/A _5299_/X vssd1 vssd1 vccd1 vccd1
+ _5388_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7127_ _7127_/CLK _7127_/D vssd1 vssd1 vccd1 vccd1 _7127_/Q sky130_fd_sc_hd__dfxtp_1
X_4339_ _4339_/A vssd1 vssd1 vccd1 vccd1 _7362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7058_ _7058_/CLK _7058_/D vssd1 vssd1 vccd1 vccd1 _7058_/Q sky130_fd_sc_hd__dfxtp_1
X_6009_ _5882_/A _6008_/X _5833_/A vssd1 vssd1 vccd1 vccd1 _6009_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6958__45 _6962__49/A vssd1 vssd1 vccd1 vccd1 _7701_/CLK sky130_fd_sc_hd__inv_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5810__299 _5810__299/A vssd1 vssd1 vccd1 vccd1 _7217_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6692__132 _6694__134/A vssd1 vssd1 vccd1 vccd1 _7576_/CLK sky130_fd_sc_hd__inv_2
X_3710_ _4095_/A _4587_/B _4039_/C vssd1 vssd1 vccd1 vccd1 _3797_/C sky130_fd_sc_hd__and3b_4
XFILLER_61_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4690_ _3813_/X _7212_/Q _4694_/S vssd1 vssd1 vccd1 vccd1 _4691_/A sky130_fd_sc_hd__mux2_1
X_3641_ _3633_/X _7690_/Q _3657_/S vssd1 vssd1 vccd1 vccd1 _3642_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3572_ _3756_/A _4376_/B _3574_/A _4376_/D vssd1 vssd1 vccd1 vccd1 _3573_/B sky130_fd_sc_hd__o22a_1
X_5311_ _5311_/A _5311_/B vssd1 vssd1 vccd1 vccd1 _5312_/A sky130_fd_sc_hd__or2_1
XFILLER_88_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5242_ _7730_/Q vssd1 vssd1 vccd1 vccd1 _6119_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_68_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5173_ _5173_/A vssd1 vssd1 vccd1 vccd1 _5360_/A sky130_fd_sc_hd__clkbuf_2
X_4124_ _4124_/A vssd1 vssd1 vccd1 vccd1 _7447_/D sky130_fd_sc_hd__clkbuf_1
X_6637__88 _6637__88/A vssd1 vssd1 vccd1 vccd1 _7532_/CLK sky130_fd_sc_hd__inv_2
Xinput1 caravel_uart_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
X_4055_ _4055_/A vssd1 vssd1 vccd1 vccd1 _7473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4957_ _5555_/B _5102_/C _5450_/A vssd1 vssd1 vccd1 vccd1 _5014_/A sky130_fd_sc_hd__and3_4
X_3908_ _3908_/A vssd1 vssd1 vccd1 vccd1 _3908_/X sky130_fd_sc_hd__buf_4
X_7676_ _7676_/CLK _7676_/D vssd1 vssd1 vccd1 vccd1 _7676_/Q sky130_fd_sc_hd__dfxtp_1
X_4888_ _4828_/X _7077_/Q _4892_/S vssd1 vssd1 vccd1 vccd1 _4889_/A sky130_fd_sc_hd__mux2_1
X_3839_ _3839_/A vssd1 vssd1 vccd1 vccd1 _7583_/D sky130_fd_sc_hd__clkbuf_1
X_6558_ _6562_/A _6558_/B _7502_/Q _6558_/D vssd1 vssd1 vccd1 vccd1 _6576_/D sky130_fd_sc_hd__and4_1
X_6489_ _7730_/Q _7499_/Q vssd1 vssd1 vccd1 vccd1 _6490_/S sky130_fd_sc_hd__xnor2_1
X_6016__303 _6017__304/A vssd1 vssd1 vccd1 vccd1 _7229_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3080_ clkbuf_0__3080_/X vssd1 vssd1 vccd1 vccd1 _6282__424/A sky130_fd_sc_hd__clkbuf_16
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2719_ clkbuf_0__2719_/X vssd1 vssd1 vccd1 vccd1 _5716__267/A sky130_fd_sc_hd__clkbuf_16
X_5860_ _5921_/A vssd1 vssd1 vccd1 vccd1 _5860_/X sky130_fd_sc_hd__clkbuf_4
X_4811_ _4811_/A vssd1 vssd1 vccd1 vccd1 _7134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5791_ _5791_/A vssd1 vssd1 vccd1 vccd1 _7204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7530_ _7530_/CLK _7530_/D vssd1 vssd1 vccd1 vccd1 _7530_/Q sky130_fd_sc_hd__dfxtp_2
X_4742_ _7165_/Q _4334_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4743_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _4673_/A vssd1 vssd1 vccd1 vccd1 _7228_/D sky130_fd_sc_hd__clkbuf_1
X_7461_ _7461_/CLK _7461_/D vssd1 vssd1 vccd1 vccd1 _7461_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__3416_ clkbuf_0__3416_/X vssd1 vssd1 vccd1 vccd1 _6937__29/A sky130_fd_sc_hd__clkbuf_16
XFILLER_119_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3624_ _3534_/X _7694_/Q _3624_/S vssd1 vssd1 vccd1 vccd1 _3625_/A sky130_fd_sc_hd__mux2_1
X_7392_ _7392_/CLK _7392_/D vssd1 vssd1 vccd1 vccd1 _7392_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__3278_ clkbuf_0__3278_/X vssd1 vssd1 vccd1 vccd1 _6685__127/A sky130_fd_sc_hd__clkbuf_16
X_6375__499 _6375__499/A vssd1 vssd1 vccd1 vccd1 _7441_/CLK sky130_fd_sc_hd__inv_2
X_3555_ _4301_/A _4561_/A _4561_/B vssd1 vssd1 vccd1 vccd1 _4882_/A sky130_fd_sc_hd__nand3_4
XFILLER_115_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3486_ _7319_/Q _7314_/Q vssd1 vssd1 vccd1 vccd1 _4467_/B sky130_fd_sc_hd__xnor2_1
X_6274_ _6274_/A _6274_/B vssd1 vssd1 vccd1 vccd1 _7359_/D sky130_fd_sc_hd__nor2_1
XFILLER_103_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5225_ _5362_/S vssd1 vssd1 vccd1 vccd1 _5225_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5156_ _7286_/Q _7072_/Q _7699_/Q _7360_/Q _5210_/A _4382_/C vssd1 vssd1 vccd1 vccd1
+ _5156_/X sky130_fd_sc_hd__mux4_1
X_5087_ _5087_/A vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__clkbuf_1
X_4107_ _4106_/X _7452_/Q _4110_/S vssd1 vssd1 vccd1 vccd1 _4108_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4038_ _4038_/A vssd1 vssd1 vccd1 vccd1 _7480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6699__138 _6700__139/A vssd1 vssd1 vccd1 vccd1 _7582_/CLK sky130_fd_sc_hd__inv_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5989_ _5882_/A _5988_/X _5833_/A vssd1 vssd1 vccd1 vccd1 _5989_/Y sky130_fd_sc_hd__o21ai_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7728_ _7731_/CLK _7728_/D vssd1 vssd1 vccd1 vccd1 _7728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7659_ _7727_/CLK _7659_/D vssd1 vssd1 vccd1 vccd1 _7659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput190 _5437_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5010_/A _5012_/B vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__and2_1
XFILLER_97_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5912_ _5912_/A vssd1 vssd1 vccd1 vccd1 _5912_/X sky130_fd_sc_hd__buf_4
X_6892_ _6903_/B vssd1 vssd1 vccd1 vccd1 _6892_/X sky130_fd_sc_hd__clkbuf_2
X_5843_ _7210_/Q _7036_/Q _7258_/Q _7250_/Q _5870_/A _5857_/A vssd1 vssd1 vccd1 vccd1
+ _5843_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5774_ _5018_/A _7197_/Q _5776_/S vssd1 vssd1 vccd1 vccd1 _5775_/A sky130_fd_sc_hd__mux2_1
X_7513_ _7525_/CLK _7513_/D vssd1 vssd1 vccd1 vccd1 _7513_/Q sky130_fd_sc_hd__dfxtp_1
X_4725_ _4725_/A vssd1 vssd1 vccd1 vccd1 _7173_/D sky130_fd_sc_hd__clkbuf_1
X_4656_ _4258_/X _7235_/Q _4658_/S vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__mux2_1
X_7444_ _7444_/CLK _7444_/D vssd1 vssd1 vccd1 vccd1 _7444_/Q sky130_fd_sc_hd__dfxtp_1
X_4587_ _4039_/C _4587_/B _4587_/C vssd1 vssd1 vccd1 vccd1 _4936_/B sky130_fd_sc_hd__and3b_2
X_3607_ _7319_/Q vssd1 vssd1 vccd1 vccd1 _4587_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput81 wbs_data_i[5] vssd1 vssd1 vccd1 vccd1 _6919_/A sky130_fd_sc_hd__buf_8
Xinput70 wbs_data_i[24] vssd1 vssd1 vccd1 vccd1 _5029_/A sky130_fd_sc_hd__buf_4
X_7375_ _7375_/CLK _7375_/D vssd1 vssd1 vccd1 vccd1 _7375_/Q sky130_fd_sc_hd__dfxtp_1
X_3538_ _3917_/A vssd1 vssd1 vccd1 vccd1 _3538_/X sky130_fd_sc_hd__buf_2
X_6326_ _6357_/A vssd1 vssd1 vccd1 vccd1 _6326_/X sky130_fd_sc_hd__buf_1
XFILLER_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3469_ _3899_/A vssd1 vssd1 vccd1 vccd1 _3469_/X sky130_fd_sc_hd__buf_2
X_5208_ _7518_/Q _5397_/S _5207_/X vssd1 vssd1 vccd1 vccd1 _5208_/X sky130_fd_sc_hd__o21ba_1
X_5139_ _5303_/A vssd1 vssd1 vccd1 vccd1 _5148_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6758__10 _6762__14/A vssd1 vssd1 vccd1 vccd1 _7629_/CLK sky130_fd_sc_hd__inv_2
X_6029__313 _6030__314/A vssd1 vssd1 vccd1 vccd1 _7239_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4510_ _7300_/Q _4325_/X _4516_/S vssd1 vssd1 vccd1 vccd1 _4511_/A sky130_fd_sc_hd__mux2_1
X_5490_ _5375_/X _7208_/Q input26/X _5376_/X vssd1 vssd1 vccd1 vccd1 _5490_/X sky130_fd_sc_hd__a22o_1
X_4441_ _4587_/C _4445_/A _6233_/A vssd1 vssd1 vccd1 vccd1 _4441_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7160_ _7160_/CLK _7160_/D vssd1 vssd1 vccd1 vccd1 _7160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4372_ _7348_/Q vssd1 vssd1 vccd1 vccd1 _5303_/A sky130_fd_sc_hd__clkbuf_2
X_6111_ _7717_/Q _7654_/Q vssd1 vssd1 vccd1 vccd1 _6792_/A sky130_fd_sc_hd__xnor2_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7723_/CLK _7091_/D vssd1 vssd1 vccd1 vccd1 _7091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6875_ _7655_/Q _6870_/X _6874_/Y vssd1 vssd1 vccd1 vccd1 _7655_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5826_ _7622_/Q _7614_/Q _7598_/Q _7590_/Q _5818_/X _5819_/X vssd1 vssd1 vccd1 vccd1
+ _5826_/X sky130_fd_sc_hd__mux4_2
XFILLER_22_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5757_ _5757_/A vssd1 vssd1 vccd1 vccd1 _7189_/D sky130_fd_sc_hd__clkbuf_1
X_4708_ _4578_/X _7180_/Q _4712_/S vssd1 vssd1 vccd1 vccd1 _4709_/A sky130_fd_sc_hd__mux2_1
X_7427_ _7427_/CLK _7427_/D vssd1 vssd1 vccd1 vccd1 _7427_/Q sky130_fd_sc_hd__dfxtp_1
X_5688_ _5688_/A vssd1 vssd1 vccd1 vccd1 _5688_/X sky130_fd_sc_hd__buf_1
X_4639_ _4639_/A vssd1 vssd1 vccd1 vccd1 _7243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7358_ _7723_/CLK _7358_/D vssd1 vssd1 vccd1 vccd1 _7358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7289_ _7289_/CLK _7289_/D vssd1 vssd1 vccd1 vccd1 _7289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__2967_ clkbuf_0__2967_/X vssd1 vssd1 vccd1 vccd1 _6175__359/A sky130_fd_sc_hd__clkbuf_16
X_6332__464 _6332__464/A vssd1 vssd1 vccd1 vccd1 _7406_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _6923_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4991_/A sky130_fd_sc_hd__and2_1
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3941_ _3660_/X _7544_/Q _3945_/S vssd1 vssd1 vccd1 vccd1 _3942_/A sky130_fd_sc_hd__mux2_1
X_3872_ _3744_/X _7569_/Q _3872_/S vssd1 vssd1 vccd1 vccd1 _3873_/A sky130_fd_sc_hd__mux2_1
X_5611_ _7089_/Q _5068_/A _5613_/S vssd1 vssd1 vccd1 vccd1 _5612_/A sky130_fd_sc_hd__mux2_1
X_6591_ _6594_/A _6592_/B vssd1 vssd1 vccd1 vccd1 _6604_/C sky130_fd_sc_hd__and2_1
X_5542_ _6913_/A _7063_/Q _5546_/S vssd1 vssd1 vccd1 vccd1 _5543_/A sky130_fd_sc_hd__mux2_1
X_5473_ _7715_/Q _5438_/X _5469_/X _5472_/X vssd1 vssd1 vccd1 vccd1 _5473_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3271_ _6645_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3271_/X sky130_fd_sc_hd__clkbuf_16
X_7212_ _7212_/CLK _7212_/D vssd1 vssd1 vccd1 vccd1 _7212_/Q sky130_fd_sc_hd__dfxtp_1
X_4424_ _4220_/X _7336_/Q _4428_/S vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__mux2_1
X_7143_ _7143_/CLK _7143_/D vssd1 vssd1 vccd1 vccd1 _7143_/Q sky130_fd_sc_hd__dfxtp_1
X_4355_ _3574_/A _4350_/B _4561_/A vssd1 vssd1 vccd1 vccd1 _4356_/C sky130_fd_sc_hd__a21o_1
XFILLER_101_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7074_ _7074_/CLK _7074_/D vssd1 vssd1 vccd1 vccd1 _7074_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _4286_/A vssd1 vssd1 vccd1 vccd1 _7383_/D sky130_fd_sc_hd__clkbuf_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6025_ _6031_/A vssd1 vssd1 vccd1 vccd1 _6025_/X sky130_fd_sc_hd__buf_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6858_ _6863_/C _6857_/C _7651_/Q vssd1 vssd1 vccd1 vccd1 _6859_/B sky130_fd_sc_hd__a21o_1
XFILLER_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6789_ _6789_/A _6789_/B _6788_/X _6135_/C vssd1 vssd1 vccd1 vccd1 _6789_/X sky130_fd_sc_hd__or4bb_1
X_6275__418 _6275__418/A vssd1 vssd1 vccd1 vccd1 _7360_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_61 _3923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_50 _3594_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_72 _7184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_83 _3549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__3097_ clkbuf_0__3097_/X vssd1 vssd1 vccd1 vccd1 _6368__493/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4140_ _4155_/S vssd1 vssd1 vccd1 vccd1 _4149_/S sky130_fd_sc_hd__buf_2
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4071_ _4071_/A vssd1 vssd1 vccd1 vccd1 _7466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4973_ _4973_/A vssd1 vssd1 vccd1 vccd1 _4973_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3924_ _3923_/X _7550_/Q _3924_/S vssd1 vssd1 vccd1 vccd1 _3925_/A sky130_fd_sc_hd__mux2_1
X_7692_ _7692_/CLK _7692_/D vssd1 vssd1 vccd1 vccd1 _7692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3855_ _3855_/A vssd1 vssd1 vccd1 vccd1 _7576_/D sky130_fd_sc_hd__clkbuf_1
X_3786_ _3744_/X _7601_/Q _3786_/S vssd1 vssd1 vccd1 vccd1 _3787_/A sky130_fd_sc_hd__mux2_1
X_6574_ _7506_/Q _6589_/B _6594_/C vssd1 vssd1 vccd1 vccd1 _6574_/X sky130_fd_sc_hd__and3_1
XFILLER_117_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5456_ _5444_/X _7189_/Q _5450_/X input5/X vssd1 vssd1 vccd1 vccd1 _5456_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XCaravelHost_195 vssd1 vssd1 vccd1 vccd1 CaravelHost_195/HI core0Index[2] sky130_fd_sc_hd__conb_1
X_4407_ _4407_/A vssd1 vssd1 vccd1 vccd1 _7344_/D sky130_fd_sc_hd__clkbuf_1
X_5387_ _5264_/X _5386_/X _4368_/A vssd1 vssd1 vccd1 vccd1 _5387_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7126_ _7126_/CLK _7126_/D vssd1 vssd1 vccd1 vccd1 _7126_/Q sky130_fd_sc_hd__dfxtp_1
X_4338_ _7362_/Q _4337_/X _4344_/S vssd1 vssd1 vccd1 vccd1 _4339_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4269_ _7390_/Q _3585_/X _4275_/S vssd1 vssd1 vccd1 vccd1 _4270_/A sky130_fd_sc_hd__mux2_1
X_7057_ _7057_/CLK _7057_/D vssd1 vssd1 vccd1 vccd1 _7057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6008_ _5929_/X _6001_/Y _6003_/Y _6005_/Y _6007_/Y vssd1 vssd1 vccd1 vccd1 _6008_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_55_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6756__9 _6756__9/A vssd1 vssd1 vccd1 vccd1 _7628_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2666_ clkbuf_0__2666_/X vssd1 vssd1 vccd1 vccd1 _5649__213/A sky130_fd_sc_hd__clkbuf_16
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6182__364 _6182__364/A vssd1 vssd1 vccd1 vccd1 _7294_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3640_ _3669_/S vssd1 vssd1 vccd1 vccd1 _3657_/S sky130_fd_sc_hd__buf_2
Xclkbuf_1_0__f__3294_ clkbuf_0__3294_/X vssd1 vssd1 vccd1 vccd1 _6925__19/A sky130_fd_sc_hd__clkbuf_16
X_3571_ _7355_/Q _7350_/Q vssd1 vssd1 vccd1 vccd1 _4376_/D sky130_fd_sc_hd__xnor2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5310_ _5281_/X _5236_/X _5308_/Y _5309_/X _5112_/X vssd1 vssd1 vccd1 vccd1 _5311_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5241_ _5375_/A _7063_/Q _5376_/A input25/X vssd1 vssd1 vccd1 vccd1 _5278_/A sky130_fd_sc_hd__a22o_1
X_5722__272 _5724__274/A vssd1 vssd1 vccd1 vccd1 _7166_/CLK sky130_fd_sc_hd__inv_2
X_5172_ _7170_/Q _7302_/Q _7488_/Q _7178_/Q _5173_/A _5171_/X vssd1 vssd1 vccd1 vccd1
+ _5172_/X sky130_fd_sc_hd__mux4_1
X_4123_ _4094_/X _7447_/Q _4131_/S vssd1 vssd1 vccd1 vccd1 _4124_/A sky130_fd_sc_hd__mux2_1
Xinput2 caravel_wb_ack_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
X_4054_ _3920_/X _7473_/Q _4056_/S vssd1 vssd1 vccd1 vccd1 _4055_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4956_ _7044_/Q _5191_/A vssd1 vssd1 vccd1 vccd1 _5450_/A sky130_fd_sc_hd__nor2_4
X_3907_ _3907_/A vssd1 vssd1 vccd1 vccd1 _7556_/D sky130_fd_sc_hd__clkbuf_1
X_7675_ _7675_/CLK _7675_/D vssd1 vssd1 vccd1 vccd1 _7675_/Q sky130_fd_sc_hd__dfxtp_1
X_4887_ _4887_/A vssd1 vssd1 vccd1 vccd1 _7078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3838_ _3750_/X _7583_/Q _3840_/S vssd1 vssd1 vccd1 vccd1 _3839_/A sky130_fd_sc_hd__mux2_1
X_6626_ _6651_/A vssd1 vssd1 vccd1 vccd1 _6626_/X sky130_fd_sc_hd__buf_1
X_6557_ _6555_/X _6556_/X _6539_/X vssd1 vssd1 vccd1 vccd1 _7503_/D sky130_fd_sc_hd__o21a_1
X_3769_ _3769_/A vssd1 vssd1 vccd1 vccd1 _7609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6488_ _7498_/Q _5235_/X vssd1 vssd1 vccd1 vccd1 _6488_/X sky130_fd_sc_hd__or2b_1
XFILLER_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5439_ _5592_/D vssd1 vssd1 vccd1 vccd1 _5493_/S sky130_fd_sc_hd__inv_2
XFILLER_105_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5578__209 _5578__209/A vssd1 vssd1 vccd1 vccd1 _7077_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7109_ _7109_/CLK _7109_/D vssd1 vssd1 vccd1 vccd1 _7109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3099_ _6376_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3099_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7722_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5665__226 _5668__229/A vssd1 vssd1 vccd1 vccd1 _7120_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2718_ clkbuf_0__2718_/X vssd1 vssd1 vccd1 vccd1 _5711__263/A sky130_fd_sc_hd__clkbuf_16
X_6642__92 _6642__92/A vssd1 vssd1 vccd1 vccd1 _7536_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4810_ _4572_/X _7134_/Q _4812_/S vssd1 vssd1 vccd1 vccd1 _4811_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5790_ _7204_/Q _5033_/A _5794_/S vssd1 vssd1 vccd1 vccd1 _5791_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4741_/A vssd1 vssd1 vccd1 vccd1 _7166_/D sky130_fd_sc_hd__clkbuf_1
X_4672_ _3813_/X _7228_/Q _4676_/S vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__mux2_1
X_7460_ _7460_/CLK _7460_/D vssd1 vssd1 vccd1 vccd1 _7460_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__3415_ clkbuf_0__3415_/X vssd1 vssd1 vccd1 vccd1 _6931__24/A sky130_fd_sc_hd__clkbuf_16
X_3623_ _3623_/A vssd1 vssd1 vccd1 vccd1 _7695_/D sky130_fd_sc_hd__clkbuf_1
X_7391_ _7391_/CLK _7391_/D vssd1 vssd1 vccd1 vccd1 _7391_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__3277_ clkbuf_0__3277_/X vssd1 vssd1 vccd1 vccd1 _6681__124/A sky130_fd_sc_hd__clkbuf_16
X_3554_ _7354_/Q vssd1 vssd1 vccd1 vccd1 _4561_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3485_ _7313_/Q vssd1 vssd1 vccd1 vccd1 _3485_/Y sky130_fd_sc_hd__clkinv_2
X_6273_ _6273_/A vssd1 vssd1 vccd1 vccd1 _7358_/D sky130_fd_sc_hd__clkbuf_1
X_5224_ _5319_/A _5224_/B vssd1 vssd1 vccd1 vccd1 _5224_/Y sky130_fd_sc_hd__nor2_1
X_5155_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5210_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5086_ _7196_/Q _5090_/B vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__and2_1
X_4106_ _7671_/Q vssd1 vssd1 vccd1 vccd1 _4106_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4037_ _3923_/X _7480_/Q _4037_/S vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _5901_/S _5981_/Y _5983_/Y _5985_/Y _5987_/Y vssd1 vssd1 vccd1 vccd1 _5988_/X
+ sky130_fd_sc_hd__o32a_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4939_ _4939_/A vssd1 vssd1 vccd1 vccd1 _7043_/D sky130_fd_sc_hd__clkbuf_1
X_7727_ _7727_/CLK _7727_/D vssd1 vssd1 vccd1 vccd1 _7727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7658_ _7731_/CLK _7658_/D vssd1 vssd1 vccd1 vccd1 _7658_/Q sky130_fd_sc_hd__dfxtp_1
X_5729__278 _5730__279/A vssd1 vssd1 vccd1 vccd1 _7172_/CLK sky130_fd_sc_hd__inv_2
X_6609_ _6609_/A _6610_/B _6609_/C vssd1 vssd1 vccd1 vccd1 _6609_/X sky130_fd_sc_hd__and3_1
X_7589_ _7589_/CLK _7589_/D vssd1 vssd1 vccd1 vccd1 _7589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_opt_1_0_wb_clk_i _7359_/CLK vssd1 vssd1 vccd1 vccd1 _6419_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput180 _5487_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput191 _5446_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6255__405 _6256__406/A vssd1 vssd1 vccd1 vccd1 _7345_/CLK sky130_fd_sc_hd__inv_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5526__196 _5529__199/A vssd1 vssd1 vccd1 vccd1 _7053_/CLK sky130_fd_sc_hd__inv_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5911_ _5906_/X _5909_/X _5995_/S vssd1 vssd1 vccd1 vccd1 _5911_/X sky130_fd_sc_hd__mux2_2
XFILLER_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6891_ _7659_/Q _6893_/B _6890_/X _6880_/X vssd1 vssd1 vccd1 vccd1 _7659_/D sky130_fd_sc_hd__o211a_1
X_5842_ _7242_/Q _7226_/Q _7472_/Q _7464_/Q _5924_/A _5841_/X vssd1 vssd1 vccd1 vccd1
+ _5842_/X sky130_fd_sc_hd__mux4_1
X_6925__19 _6925__19/A vssd1 vssd1 vccd1 vccd1 _7675_/CLK sky130_fd_sc_hd__inv_2
X_5773_ _5773_/A vssd1 vssd1 vccd1 vccd1 _7196_/D sky130_fd_sc_hd__clkbuf_1
X_4724_ _4575_/X _7173_/Q _4724_/S vssd1 vssd1 vccd1 vccd1 _4725_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7512_ _7525_/CLK _7512_/D vssd1 vssd1 vccd1 vccd1 _7512_/Q sky130_fd_sc_hd__dfxtp_1
X_4655_ _4655_/A vssd1 vssd1 vccd1 vccd1 _7236_/D sky130_fd_sc_hd__clkbuf_1
X_7443_ _7443_/CLK _7443_/D vssd1 vssd1 vccd1 vccd1 _7443_/Q sky130_fd_sc_hd__dfxtp_1
X_3606_ _3900_/C vssd1 vssd1 vccd1 vccd1 _4039_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4586_ _4586_/A vssd1 vssd1 vccd1 vccd1 _7266_/D sky130_fd_sc_hd__clkbuf_1
Xinput82 wbs_data_i[6] vssd1 vssd1 vccd1 vccd1 _6921_/A sky130_fd_sc_hd__buf_8
Xinput60 wbs_data_i[15] vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__buf_4
Xinput71 wbs_data_i[25] vssd1 vssd1 vccd1 vccd1 _5031_/A sky130_fd_sc_hd__buf_4
X_7374_ _7374_/CLK _7374_/D vssd1 vssd1 vccd1 vccd1 _7374_/Q sky130_fd_sc_hd__dfxtp_1
X_3537_ _7669_/Q vssd1 vssd1 vccd1 vccd1 _3917_/A sky130_fd_sc_hd__buf_2
X_3468_ _7674_/Q vssd1 vssd1 vccd1 vccd1 _3899_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5207_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__buf_2
XFILLER_57_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5138_ _5429_/S vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5069_ _5069_/A vssd1 vssd1 vccd1 vccd1 _5069_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4440_ _4587_/B _4443_/A _4443_/B vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__and3_1
X_6110_ _6458_/B vssd1 vssd1 vccd1 vccd1 _6112_/A sky130_fd_sc_hd__clkbuf_2
X_4371_ _5415_/A vssd1 vssd1 vccd1 vccd1 _5315_/A sky130_fd_sc_hd__clkbuf_2
X_7090_ _7190_/CLK _7090_/D vssd1 vssd1 vccd1 vccd1 _7090_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5678__236 _5681__239/A vssd1 vssd1 vccd1 vccd1 _7130_/CLK sky130_fd_sc_hd__inv_2
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6874_ _7655_/Q _6870_/X _6864_/A vssd1 vssd1 vccd1 vccd1 _6874_/Y sky130_fd_sc_hd__a21oi_1
X_5825_ _5899_/S _5825_/B vssd1 vssd1 vccd1 vccd1 _5825_/X sky130_fd_sc_hd__or2_1
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5756_ _4999_/A _7189_/Q _5758_/S vssd1 vssd1 vccd1 vccd1 _5757_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4707_ _4707_/A vssd1 vssd1 vccd1 vccd1 _7181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4638_ _4258_/X _7243_/Q _4640_/S vssd1 vssd1 vccd1 vccd1 _4639_/A sky130_fd_sc_hd__mux2_1
X_7426_ _7426_/CLK _7426_/D vssd1 vssd1 vccd1 vccd1 _7426_/Q sky130_fd_sc_hd__dfxtp_1
X_6203__381 _6204__382/A vssd1 vssd1 vccd1 vccd1 _7311_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4569_ _4569_/A vssd1 vssd1 vccd1 vccd1 _4569_/X sky130_fd_sc_hd__clkbuf_4
X_7357_ _7357_/CLK _7357_/D vssd1 vssd1 vccd1 vccd1 _7357_/Q sky130_fd_sc_hd__dfxtp_1
X_6308_ _6308_/A vssd1 vssd1 vccd1 vccd1 _6308_/X sky130_fd_sc_hd__buf_1
X_7288_ _7288_/CLK _7288_/D vssd1 vssd1 vccd1 vccd1 _7288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2966_ clkbuf_0__2966_/X vssd1 vssd1 vccd1 vccd1 _6083__352/A sky130_fd_sc_hd__clkbuf_16
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6408__525 _6412__529/A vssd1 vssd1 vccd1 vccd1 _7467_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3940_ _3940_/A vssd1 vssd1 vccd1 vccd1 _7545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3871_ _3871_/A vssd1 vssd1 vccd1 vccd1 _7570_/D sky130_fd_sc_hd__clkbuf_1
X_6656__104 _6656__104/A vssd1 vssd1 vccd1 vccd1 _7548_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5610_ _5610_/A vssd1 vssd1 vccd1 vccd1 _7088_/D sky130_fd_sc_hd__clkbuf_1
X_6590_ _6588_/X _6589_/X _6569_/X vssd1 vssd1 vccd1 vccd1 _7509_/D sky130_fd_sc_hd__o21a_1
X_5541_ _5541_/A vssd1 vssd1 vccd1 vccd1 _7062_/D sky130_fd_sc_hd__clkbuf_1
X_7211_ _7211_/CLK _7211_/D vssd1 vssd1 vccd1 vccd1 _7211_/Q sky130_fd_sc_hd__dfxtp_1
X_5472_ _5375_/A _7195_/Q input11/X _5102_/D vssd1 vssd1 vccd1 vccd1 _5472_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_0__3270_ _6639_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3270_/X sky130_fd_sc_hd__clkbuf_16
X_4423_ _4423_/A vssd1 vssd1 vccd1 vccd1 _7337_/D sky130_fd_sc_hd__clkbuf_1
X_4354_ _6222_/A vssd1 vssd1 vccd1 vccd1 _6272_/C sky130_fd_sc_hd__clkbuf_2
X_7142_ _7142_/CLK _7142_/D vssd1 vssd1 vccd1 vccd1 _7142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7073_ _7073_/CLK _7073_/D vssd1 vssd1 vccd1 vccd1 _7073_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _6055_/A vssd1 vssd1 vccd1 vccd1 _6024_/X sky130_fd_sc_hd__buf_1
X_4285_ _4238_/X _7383_/Q _4293_/S vssd1 vssd1 vccd1 vccd1 _4286_/A sky130_fd_sc_hd__mux2_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _6932_/A vssd1 vssd1 vccd1 vccd1 _6926_/X sky130_fd_sc_hd__buf_1
XFILLER_82_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6309__445 _6313__449/A vssd1 vssd1 vccd1 vccd1 _7387_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6857_ _7651_/Q _6863_/C _6857_/C vssd1 vssd1 vccd1 vccd1 _6857_/X sky130_fd_sc_hd__and3_1
XFILLER_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6788_ _6788_/A _6788_/B _6788_/C vssd1 vssd1 vccd1 vccd1 _6788_/X sky130_fd_sc_hd__and3_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5739_ _5745_/A vssd1 vssd1 vccd1 vccd1 _5739_/X sky130_fd_sc_hd__buf_1
XFILLER_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7409_ _7409_/CLK _7409_/D vssd1 vssd1 vccd1 vccd1 _7409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_51 _3603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_40 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_84 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_73 _7543_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_62 _4331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3096_ clkbuf_0__3096_/X vssd1 vssd1 vccd1 vccd1 _6363__489/A sky130_fd_sc_hd__clkbuf_16
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6649__98 _6650__99/A vssd1 vssd1 vccd1 vccd1 _7542_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _3917_/X _7466_/Q _4074_/S vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6380__503 _6381__504/A vssd1 vssd1 vccd1 vccd1 _7445_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4972_ _5784_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4973_/A sky130_fd_sc_hd__and2_1
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3923_ _3923_/A vssd1 vssd1 vccd1 vccd1 _3923_/X sky130_fd_sc_hd__buf_4
X_7691_ _7691_/CLK _7691_/D vssd1 vssd1 vccd1 vccd1 _7691_/Q sky130_fd_sc_hd__dfxtp_1
X_3854_ _3747_/X _7576_/Q _3858_/S vssd1 vssd1 vccd1 vccd1 _3855_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3785_ _3785_/A vssd1 vssd1 vccd1 vccd1 _7602_/D sky130_fd_sc_hd__clkbuf_1
X_6573_ _6571_/A _6571_/B _6577_/B _6607_/B _6609_/C vssd1 vssd1 vccd1 vccd1 _6573_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_118_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5524_ _5573_/A vssd1 vssd1 vccd1 vccd1 _5524_/X sky130_fd_sc_hd__buf_1
X_5455_ _6129_/A _5448_/X _5449_/X _5454_/X vssd1 vssd1 vccd1 vccd1 _5455_/X sky130_fd_sc_hd__a31o_1
XCaravelHost_196 vssd1 vssd1 vccd1 vccd1 CaravelHost_196/HI core0Index[3] sky130_fd_sc_hd__conb_1
X_4406_ _7344_/Q _4328_/X _4410_/S vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7125_ _7125_/CLK _7125_/D vssd1 vssd1 vccd1 vccd1 _7125_/Q sky130_fd_sc_hd__dfxtp_1
X_5386_ _7374_/Q _7345_/Q _7337_/Q _7300_/Q _5290_/S _5365_/A vssd1 vssd1 vccd1 vccd1
+ _5386_/X sky130_fd_sc_hd__mux4_1
X_4337_ _7323_/Q vssd1 vssd1 vccd1 vccd1 _4337_/X sky130_fd_sc_hd__buf_4
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7056_ _7056_/CLK _7056_/D vssd1 vssd1 vccd1 vccd1 _7056_/Q sky130_fd_sc_hd__dfxtp_1
X_4268_ _4268_/A vssd1 vssd1 vccd1 vccd1 _7391_/D sky130_fd_sc_hd__clkbuf_1
X_6007_ _5923_/A _6006_/X _5917_/A vssd1 vssd1 vccd1 vccd1 _6007_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4199_ _4103_/X _7413_/Q _4203_/S vssd1 vssd1 vccd1 vccd1 _4200_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6281__423 _6281__423/A vssd1 vssd1 vccd1 vccd1 _7365_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6909_/A vssd1 vssd1 vccd1 vccd1 _7667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__2665_ clkbuf_0__2665_/X vssd1 vssd1 vccd1 vccd1 _5669_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3293_ clkbuf_0__3293_/X vssd1 vssd1 vccd1 vccd1 _6762__14/A sky130_fd_sc_hd__clkbuf_16
X_3570_ _7354_/Q _7353_/Q _3570_/C vssd1 vssd1 vccd1 vccd1 _3574_/A sky130_fd_sc_hd__and3_1
XFILLER_115_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5240_ _5240_/A vssd1 vssd1 vccd1 vccd1 _5240_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5171_ _5325_/S vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__buf_2
XFILLER_110_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4137_/S vssd1 vssd1 vccd1 vccd1 _4131_/S sky130_fd_sc_hd__buf_2
X_4053_ _4053_/A vssd1 vssd1 vccd1 vccd1 _7474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 caravel_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_4
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4955_ _5591_/B vssd1 vssd1 vccd1 vccd1 _5191_/A sky130_fd_sc_hd__inv_2
X_3906_ _3905_/X _7556_/Q _3915_/S vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__mux2_1
X_7674_ _7674_/CLK _7674_/D vssd1 vssd1 vccd1 vccd1 _7674_/Q sky130_fd_sc_hd__dfxtp_1
X_4886_ _4825_/X _7078_/Q _4892_/S vssd1 vssd1 vccd1 vccd1 _4887_/A sky130_fd_sc_hd__mux2_1
X_3837_ _3837_/A vssd1 vssd1 vccd1 vccd1 _7584_/D sky130_fd_sc_hd__clkbuf_1
X_6625_ _6719_/A vssd1 vssd1 vccd1 vccd1 _6625_/X sky130_fd_sc_hd__buf_1
X_3768_ _3656_/X _7609_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3769_/A sky130_fd_sc_hd__mux2_1
X_6556_ _6558_/B _6556_/B _6562_/C vssd1 vssd1 vccd1 vccd1 _6556_/X sky130_fd_sc_hd__and3_1
X_6669__114 _6669__114/A vssd1 vssd1 vccd1 vccd1 _7558_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3699_ _3530_/X _7634_/Q _3701_/S vssd1 vssd1 vccd1 vccd1 _3700_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6487_ _6487_/A _7498_/Q vssd1 vssd1 vccd1 vccd1 _6487_/X sky130_fd_sc_hd__or2b_1
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5438_ _5494_/S vssd1 vssd1 vccd1 vccd1 _5438_/X sky130_fd_sc_hd__clkbuf_2
X_5369_ _5158_/X _5356_/Y _5361_/X _5368_/X _5161_/A vssd1 vssd1 vccd1 vccd1 _5369_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_113_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6387__509 _6387__509/A vssd1 vssd1 vccd1 vccd1 _7451_/CLK sky130_fd_sc_hd__inv_2
X_7108_ _7108_/CLK _7108_/D vssd1 vssd1 vccd1 vccd1 _7108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7039_ _7039_/CLK _7039_/D vssd1 vssd1 vccd1 vccd1 _7039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3098_ _6370_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3098_/X sky130_fd_sc_hd__clkbuf_16
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023__309 _6023__309/A vssd1 vssd1 vccd1 vccd1 _7235_/CLK sky130_fd_sc_hd__inv_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6288__429 _6288__429/A vssd1 vssd1 vccd1 vccd1 _7371_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2717_ clkbuf_0__2717_/X vssd1 vssd1 vccd1 vccd1 _5731_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_19_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4740_ _7166_/Q _4331_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4741_/A sky130_fd_sc_hd__mux2_1
X_4671_ _4671_/A vssd1 vssd1 vccd1 vccd1 _7229_/D sky130_fd_sc_hd__clkbuf_1
X_3622_ _3530_/X _7695_/Q _3624_/S vssd1 vssd1 vccd1 vccd1 _3623_/A sky130_fd_sc_hd__mux2_1
X_7390_ _7390_/CLK _7390_/D vssd1 vssd1 vccd1 vccd1 _7390_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__3276_ clkbuf_0__3276_/X vssd1 vssd1 vccd1 vccd1 _6674__118/A sky130_fd_sc_hd__clkbuf_16
XFILLER_115_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3553_ _3926_/A vssd1 vssd1 vccd1 vccd1 _4561_/A sky130_fd_sc_hd__buf_2
XFILLER_103_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3484_ _3484_/A _3484_/B vssd1 vssd1 vccd1 vccd1 _3494_/B sky130_fd_sc_hd__or2_1
X_6272_ _7715_/Q _7285_/Q _6272_/C vssd1 vssd1 vccd1 vccd1 _6273_/A sky130_fd_sc_hd__and3_1
X_5223_ _7543_/Q _7433_/Q _7401_/Q _7385_/Q _5330_/S _4375_/A vssd1 vssd1 vccd1 vccd1
+ _5224_/B sky130_fd_sc_hd__mux4_1
XFILLER_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5154_ _7348_/Q vssd1 vssd1 vccd1 vccd1 _5207_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4105_ _4105_/A vssd1 vssd1 vccd1 vccd1 _7453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5085_ _5085_/A vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4036_ _4036_/A vssd1 vssd1 vccd1 vccd1 _7481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5987_ _5923_/A _5986_/X _5929_/X vssd1 vssd1 vccd1 vccd1 _5987_/Y sky130_fd_sc_hd__o21ai_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4938_ _3794_/X _7043_/Q _4946_/S vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__mux2_1
X_7726_ _7731_/CLK _7726_/D vssd1 vssd1 vccd1 vccd1 _7726_/Q sky130_fd_sc_hd__dfxtp_1
X_7657_ _7722_/CLK _7657_/D vssd1 vssd1 vccd1 vccd1 _7657_/Q sky130_fd_sc_hd__dfxtp_1
X_4869_ _4869_/A vssd1 vssd1 vccd1 vccd1 _7112_/D sky130_fd_sc_hd__clkbuf_1
X_6393__513 _6394__514/A vssd1 vssd1 vccd1 vccd1 _7455_/CLK sky130_fd_sc_hd__inv_2
X_6608_ _7513_/Q _6605_/Y _6606_/X _6615_/A vssd1 vssd1 vccd1 vccd1 _7513_/D sky130_fd_sc_hd__o211a_1
X_7588_ _7588_/CLK _7588_/D vssd1 vssd1 vccd1 vccd1 _7588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6539_ _6569_/A vssd1 vssd1 vccd1 vccd1 _6539_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput170 _5476_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput192 _5452_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[9] sky130_fd_sc_hd__buf_2
Xoutput181 _5488_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[28] sky130_fd_sc_hd__buf_2
XFILLER_101_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5671__231 _5673__233/A vssd1 vssd1 vccd1 vccd1 _7125_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5910_ _5910_/A vssd1 vssd1 vccd1 vccd1 _5995_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_53_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6890_ _7660_/Q _6903_/B vssd1 vssd1 vccd1 vccd1 _6890_/X sky130_fd_sc_hd__or2_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5841_ _5856_/A vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5772_ _5016_/A _7196_/Q _5776_/S vssd1 vssd1 vccd1 vccd1 _5773_/A sky130_fd_sc_hd__mux2_1
X_6739__170 _6741__172/A vssd1 vssd1 vccd1 vccd1 _7614_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4723_ _4723_/A vssd1 vssd1 vccd1 vccd1 _7174_/D sky130_fd_sc_hd__clkbuf_1
X_7511_ _7525_/CLK _7511_/D vssd1 vssd1 vccd1 vccd1 _7511_/Q sky130_fd_sc_hd__dfxtp_1
X_7442_ _7442_/CLK _7442_/D vssd1 vssd1 vccd1 vccd1 _7442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4654_ _4255_/X _7236_/Q _4658_/S vssd1 vssd1 vccd1 vccd1 _4655_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3605_ _3605_/A vssd1 vssd1 vccd1 vccd1 _7699_/D sky130_fd_sc_hd__clkbuf_1
X_4585_ _4584_/X _7266_/Q _4585_/S vssd1 vssd1 vccd1 vccd1 _4586_/A sky130_fd_sc_hd__mux2_1
Xinput50 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _5062_/A sky130_fd_sc_hd__buf_4
Xinput61 wbs_data_i[16] vssd1 vssd1 vccd1 vccd1 _5010_/A sky130_fd_sc_hd__buf_4
Xinput72 wbs_data_i[26] vssd1 vssd1 vccd1 vccd1 _5033_/A sky130_fd_sc_hd__buf_4
X_7373_ _7373_/CLK _7373_/D vssd1 vssd1 vccd1 vccd1 _7373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3536_ _3536_/A vssd1 vssd1 vccd1 vccd1 _7710_/D sky130_fd_sc_hd__clkbuf_1
Xinput83 wbs_data_i[7] vssd1 vssd1 vccd1 vccd1 _6923_/A sky130_fd_sc_hd__buf_8
XFILLER_89_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5206_ _5201_/X _5203_/X _5204_/X _5257_/A _5205_/X vssd1 vssd1 vccd1 vccd1 _5217_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5137_ _5245_/A vssd1 vssd1 vccd1 vccd1 _5429_/S sky130_fd_sc_hd__clkbuf_2
X_5068_ _5068_/A _5068_/B vssd1 vssd1 vccd1 vccd1 _5069_/A sky130_fd_sc_hd__and2_1
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4019_ _7488_/Q _3603_/X _4019_/S vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5735__283 _5735__283/A vssd1 vssd1 vccd1 vccd1 _7177_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7709_ _7709_/CLK _7709_/D vssd1 vssd1 vccd1 vccd1 _7709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2719_ _5713_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2719_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5742__287 _5744__289/A vssd1 vssd1 vccd1 vccd1 _7181_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2630_ clkbuf_0__2630_/X vssd1 vssd1 vccd1 vccd1 _5517__189/A sky130_fd_sc_hd__clkbuf_16
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6930__23 _6930__23/A vssd1 vssd1 vccd1 vccd1 _7679_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4370_ _5262_/A vssd1 vssd1 vccd1 vccd1 _5415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6036__319 _6036__319/A vssd1 vssd1 vccd1 vccd1 _7245_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6873_ _6873_/A vssd1 vssd1 vccd1 vccd1 _7654_/D sky130_fd_sc_hd__clkbuf_1
X_5824_ _7392_/Q _7234_/Q _7550_/Q _7456_/Q _5908_/A _5823_/X vssd1 vssd1 vccd1 vccd1
+ _5825_/B sky130_fd_sc_hd__mux4_1
X_6764__15 _6925__19/A vssd1 vssd1 vccd1 vccd1 _7634_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5755_ _5755_/A vssd1 vssd1 vccd1 vccd1 _7188_/D sky130_fd_sc_hd__clkbuf_1
X_4706_ _4575_/X _7181_/Q _4706_/S vssd1 vssd1 vccd1 vccd1 _4707_/A sky130_fd_sc_hd__mux2_1
X_4637_ _4637_/A vssd1 vssd1 vccd1 vccd1 _7244_/D sky130_fd_sc_hd__clkbuf_1
X_7425_ _7425_/CLK _7425_/D vssd1 vssd1 vccd1 vccd1 _7425_/Q sky130_fd_sc_hd__dfxtp_1
X_5806__295 _5810__299/A vssd1 vssd1 vccd1 vccd1 _7213_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4568_ _4568_/A vssd1 vssd1 vccd1 vccd1 _7272_/D sky130_fd_sc_hd__clkbuf_1
X_7356_ _7356_/CLK _7356_/D vssd1 vssd1 vccd1 vccd1 _7356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3519_ _3469_/X _7714_/Q _3535_/S vssd1 vssd1 vccd1 vccd1 _3520_/A sky130_fd_sc_hd__mux2_1
X_7287_ _7287_/CLK _7287_/D vssd1 vssd1 vccd1 vccd1 _7287_/Q sky130_fd_sc_hd__dfxtp_1
X_4499_ _4499_/A vssd1 vssd1 vccd1 vccd1 _7305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6889_/A _6768_/A vssd1 vssd1 vccd1 vccd1 _6805_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6210__386 _6210__386/A vssd1 vssd1 vccd1 vccd1 _7316_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3870_ _3741_/X _7570_/Q _3872_/S vssd1 vssd1 vccd1 vccd1 _3871_/A sky130_fd_sc_hd__mux2_1
X_6081__350 _6085__354/A vssd1 vssd1 vccd1 vccd1 _7279_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5540_ _6911_/A _7062_/Q _5546_/S vssd1 vssd1 vccd1 vccd1 _5541_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5684__241 _5687__244/A vssd1 vssd1 vccd1 vccd1 _7135_/CLK sky130_fd_sc_hd__inv_2
X_5471_ _7716_/Q _5438_/X _5469_/X _5470_/X vssd1 vssd1 vccd1 vccd1 _5471_/X sky130_fd_sc_hd__a31o_1
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7210_ _7210_/CLK _7210_/D vssd1 vssd1 vccd1 vccd1 _7210_/Q sky130_fd_sc_hd__dfxtp_1
X_4422_ _4217_/X _7337_/Q _4428_/S vssd1 vssd1 vccd1 vccd1 _4423_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7141_ _7141_/CLK _7141_/D vssd1 vssd1 vccd1 vccd1 _7141_/Q sky130_fd_sc_hd__dfxtp_1
X_4353_ _4301_/A _6220_/B _4356_/B _4774_/S vssd1 vssd1 vccd1 vccd1 _7356_/D sky130_fd_sc_hd__a31o_1
X_4284_ _4299_/S vssd1 vssd1 vccd1 vccd1 _4293_/S sky130_fd_sc_hd__buf_2
X_7072_ _7072_/CLK _7072_/D vssd1 vssd1 vccd1 vccd1 _7072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6663__109 _6663__109/A vssd1 vssd1 vccd1 vccd1 _7553_/CLK sky130_fd_sc_hd__inv_2
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6856_ _6856_/A vssd1 vssd1 vccd1 vccd1 _7650_/D sky130_fd_sc_hd__clkbuf_1
X_3999_ _3999_/A vssd1 vssd1 vccd1 vccd1 _7518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6787_ _6098_/Y _7650_/Q _6118_/A _5281_/X vssd1 vssd1 vccd1 vccd1 _6788_/C sky130_fd_sc_hd__o2bb2a_1
XFILLER_13_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5738_ _6207_/A vssd1 vssd1 vccd1 vccd1 _5738_/X sky130_fd_sc_hd__buf_1
XFILLER_89_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5669_ _5669_/A vssd1 vssd1 vccd1 vccd1 _5669_/X sky130_fd_sc_hd__buf_1
X_7408_ _7408_/CLK _7408_/D vssd1 vssd1 vccd1 vccd1 _7408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7339_ _7339_/CLK _7339_/D vssd1 vssd1 vccd1 vccd1 _7339_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_30 _5049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_41 _6919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_52 _6915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6425__58 _6426__59/A vssd1 vssd1 vccd1 vccd1 _7480_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_85 _3801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_74 _7545_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_63 _5481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__3095_ clkbuf_0__3095_/X vssd1 vssd1 vccd1 vccd1 _6382_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_119_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6414__530 _6416__532/A vssd1 vssd1 vccd1 vccd1 _7472_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4971_ _4971_/A vssd1 vssd1 vccd1 vccd1 _4971_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3922_ _3922_/A vssd1 vssd1 vccd1 vccd1 _7551_/D sky130_fd_sc_hd__clkbuf_1
X_7690_ _7690_/CLK _7690_/D vssd1 vssd1 vccd1 vccd1 _7690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3853_ _3853_/A vssd1 vssd1 vccd1 vccd1 _7577_/D sky130_fd_sc_hd__clkbuf_1
X_3784_ _3741_/X _7602_/Q _3786_/S vssd1 vssd1 vccd1 vccd1 _3785_/A sky130_fd_sc_hd__mux2_1
X_6572_ _6572_/A _6572_/B _6572_/C vssd1 vssd1 vccd1 vccd1 _6609_/C sky130_fd_sc_hd__and3_1
XFILLER_118_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5454_ _5444_/X _7188_/Q _5450_/X input4/X vssd1 vssd1 vccd1 vccd1 _5454_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_197 vssd1 vssd1 vccd1 vccd1 CaravelHost_197/HI core0Index[4] sky130_fd_sc_hd__conb_1
X_4405_ _4405_/A vssd1 vssd1 vccd1 vccd1 _7345_/D sky130_fd_sc_hd__clkbuf_1
X_5385_ _5291_/A _5382_/X _5384_/X _5351_/A vssd1 vssd1 vccd1 vccd1 _5385_/X sky130_fd_sc_hd__a211o_1
X_7124_ _7124_/CLK _7124_/D vssd1 vssd1 vccd1 vccd1 _7124_/Q sky130_fd_sc_hd__dfxtp_1
X_4336_ _4336_/A vssd1 vssd1 vccd1 vccd1 _7363_/D sky130_fd_sc_hd__clkbuf_1
X_6315__450 _6317__452/A vssd1 vssd1 vccd1 vccd1 _7392_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7055_ _7055_/CLK _7055_/D vssd1 vssd1 vccd1 vccd1 _7055_/Q sky130_fd_sc_hd__dfxtp_1
X_4267_ _7391_/Q _3549_/X _4275_/S vssd1 vssd1 vccd1 vccd1 _4268_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6006_ _7415_/Q _7383_/Q _7714_/Q _7637_/Q _5921_/X _5884_/X vssd1 vssd1 vccd1 vccd1
+ _6006_/X sky130_fd_sc_hd__mux4_1
X_4198_ _4198_/A vssd1 vssd1 vccd1 vccd1 _7414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6908_ _6908_/A _6923_/B vssd1 vssd1 vccd1 vccd1 _6909_/A sky130_fd_sc_hd__and2_1
Xclkbuf_0__2967_ _6086_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2967_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6839_ _6847_/C _6843_/C vssd1 vssd1 vccd1 vccd1 _6841_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2664_ clkbuf_0__2664_/X vssd1 vssd1 vccd1 vccd1 _5576__207/A sky130_fd_sc_hd__clkbuf_16
XFILLER_18_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5531__200 _5572__204/A vssd1 vssd1 vccd1 vccd1 _7057_/CLK sky130_fd_sc_hd__inv_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3292_ clkbuf_0__3292_/X vssd1 vssd1 vccd1 vccd1 _6756__9/A sky130_fd_sc_hd__clkbuf_16
X_6733__165 _6737__169/A vssd1 vssd1 vccd1 vccd1 _7609_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__3078_ clkbuf_0__3078_/X vssd1 vssd1 vccd1 vccd1 _6275__418/A sky130_fd_sc_hd__clkbuf_16
XFILLER_115_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5170_ _5270_/A vssd1 vssd1 vccd1 vccd1 _5325_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_96_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4121_ _4121_/A _4175_/B vssd1 vssd1 vccd1 vccd1 _4137_/S sky130_fd_sc_hd__or2_4
XFILLER_110_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4052_ _3917_/X _7474_/Q _4056_/S vssd1 vssd1 vccd1 vccd1 _4053_/A sky130_fd_sc_hd__mux2_1
Xinput4 caravel_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4954_ _7209_/Q _7208_/Q _7207_/Q _7206_/Q vssd1 vssd1 vccd1 vccd1 _5102_/C sky130_fd_sc_hd__and4bb_4
X_3905_ _3905_/A vssd1 vssd1 vccd1 vccd1 _3905_/X sky130_fd_sc_hd__buf_4
X_7673_ _7674_/CLK _7673_/D vssd1 vssd1 vccd1 vccd1 _7673_/Q sky130_fd_sc_hd__dfxtp_2
X_4885_ _4885_/A vssd1 vssd1 vccd1 vccd1 _7079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3836_ _3747_/X _7584_/Q _3840_/S vssd1 vssd1 vccd1 vccd1 _3837_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3767_ _3767_/A vssd1 vssd1 vccd1 vccd1 _7610_/D sky130_fd_sc_hd__clkbuf_1
X_6555_ _6559_/B _6583_/C _6555_/C vssd1 vssd1 vccd1 vccd1 _6555_/X sky130_fd_sc_hd__and3b_1
X_5506_ _5518_/A vssd1 vssd1 vccd1 vccd1 _5506_/X sky130_fd_sc_hd__buf_1
XFILLER_118_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3698_ _3698_/A vssd1 vssd1 vccd1 vccd1 _7635_/D sky130_fd_sc_hd__clkbuf_1
X_6486_ _7500_/Q _6486_/B _6486_/C vssd1 vssd1 vccd1 vccd1 _6486_/Y sky130_fd_sc_hd__nand3b_1
X_6239__392 _6240__393/A vssd1 vssd1 vccd1 vccd1 _7332_/CLK sky130_fd_sc_hd__inv_2
X_5437_ _5481_/A _7068_/Q _5482_/A input32/X _5436_/X vssd1 vssd1 vccd1 vccd1 _5437_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5368_ _5264_/X _5363_/Y _5365_/X _5367_/Y vssd1 vssd1 vccd1 vccd1 _5368_/X sky130_fd_sc_hd__a31o_1
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5299_ _5299_/A vssd1 vssd1 vccd1 vccd1 _5299_/X sky130_fd_sc_hd__clkbuf_4
X_7107_ _7107_/CLK _7107_/D vssd1 vssd1 vccd1 vccd1 _7107_/Q sky130_fd_sc_hd__dfxtp_1
X_4319_ _4319_/A vssd1 vssd1 vccd1 vccd1 _7368_/D sky130_fd_sc_hd__clkbuf_1
X_7038_ _7038_/CLK _7038_/D vssd1 vssd1 vccd1 vccd1 _7038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3097_ _6364_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3097_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6627__80 _6628__81/A vssd1 vssd1 vccd1 vccd1 _7523_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__2716_ clkbuf_0__2716_/X vssd1 vssd1 vccd1 vccd1 _5702__256/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6937__29 _6937__29/A vssd1 vssd1 vccd1 vccd1 _7685_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _3810_/X _7229_/Q _4670_/S vssd1 vssd1 vccd1 vccd1 _4671_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3621_ _3621_/A vssd1 vssd1 vccd1 vccd1 _7696_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__3275_ clkbuf_0__3275_/X vssd1 vssd1 vccd1 vccd1 _6669__114/A sky130_fd_sc_hd__clkbuf_16
X_3552_ _7355_/Q vssd1 vssd1 vccd1 vccd1 _3926_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3483_ _4443_/A _3483_/B vssd1 vssd1 vccd1 vccd1 _3494_/A sky130_fd_sc_hd__or2_1
XFILLER_102_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5222_ _5429_/S vssd1 vssd1 vccd1 vccd1 _5330_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_102_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5153_ _5163_/A vssd1 vssd1 vccd1 vccd1 _5319_/A sky130_fd_sc_hd__clkbuf_2
X_4104_ _4103_/X _7453_/Q _4110_/S vssd1 vssd1 vccd1 vccd1 _4105_/A sky130_fd_sc_hd__mux2_1
X_5084_ _7195_/Q _5090_/B vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__and2_1
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4035_ _3920_/X _7481_/Q _4037_/S vssd1 vssd1 vccd1 vccd1 _4036_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5986_ _7414_/Q _7382_/Q _7713_/Q _7636_/Q _5921_/X _5884_/X vssd1 vssd1 vccd1 vccd1
+ _5986_/X sky130_fd_sc_hd__mux4_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ _4952_/S vssd1 vssd1 vccd1 vccd1 _4946_/S sky130_fd_sc_hd__clkbuf_4
X_7725_ _7731_/CLK _7725_/D vssd1 vssd1 vccd1 vccd1 _7725_/Q sky130_fd_sc_hd__dfxtp_1
X_7656_ _7731_/CLK _7656_/D vssd1 vssd1 vccd1 vccd1 _7656_/Q sky130_fd_sc_hd__dfxtp_1
X_4868_ _4825_/X _7112_/Q _4874_/S vssd1 vssd1 vccd1 vccd1 _4869_/A sky130_fd_sc_hd__mux2_1
X_3819_ _7667_/Q vssd1 vssd1 vccd1 vccd1 _3819_/X sky130_fd_sc_hd__buf_6
X_6607_ _6607_/A _6607_/B vssd1 vssd1 vccd1 vccd1 _6615_/A sky130_fd_sc_hd__nor2_2
Xclkbuf_0__2666_ _5580_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2666_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7587_ _7587_/CLK _7587_/D vssd1 vssd1 vccd1 vccd1 _7587_/Q sky130_fd_sc_hd__dfxtp_1
X_4799_ _4799_/A vssd1 vssd1 vccd1 vccd1 _7139_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6538_ _6541_/B _6556_/B _6562_/C vssd1 vssd1 vccd1 vccd1 _6538_/X sky130_fd_sc_hd__and3_1
XFILLER_118_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6469_ _6777_/A _6470_/C _6571_/A vssd1 vssd1 vccd1 vccd1 _6469_/X sky130_fd_sc_hd__a21o_1
Xoutput160 _5495_/X vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
Xoutput182 _5489_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[29] sky130_fd_sc_hd__buf_2
Xoutput171 _5477_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[19] sky130_fd_sc_hd__buf_2
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6328__460 _6331__463/A vssd1 vssd1 vccd1 vccd1 _7402_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6942__32 _6944__34/A vssd1 vssd1 vccd1 vccd1 _7688_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6294__434 _6294__434/A vssd1 vssd1 vccd1 vccd1 _7376_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5840_ _5837_/X _5838_/X _5910_/A vssd1 vssd1 vccd1 vccd1 _5840_/X sky130_fd_sc_hd__mux2_2
X_5771_ _5771_/A vssd1 vssd1 vccd1 vccd1 _7195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4722_ _4572_/X _7174_/Q _4724_/S vssd1 vssd1 vccd1 vccd1 _4723_/A sky130_fd_sc_hd__mux2_1
X_7510_ _7510_/CLK _7510_/D vssd1 vssd1 vccd1 vccd1 _7510_/Q sky130_fd_sc_hd__dfxtp_1
X_7441_ _7441_/CLK _7441_/D vssd1 vssd1 vccd1 vccd1 _7441_/Q sky130_fd_sc_hd__dfxtp_1
X_5648__212 _5649__213/A vssd1 vssd1 vccd1 vccd1 _7106_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4653_ _4653_/A vssd1 vssd1 vccd1 vccd1 _7237_/D sky130_fd_sc_hd__clkbuf_1
Xinput40 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__buf_4
XFILLER_30_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3604_ _7699_/Q _3603_/X _3604_/S vssd1 vssd1 vccd1 vccd1 _3605_/A sky130_fd_sc_hd__mux2_1
X_4584_ _4584_/A vssd1 vssd1 vccd1 vccd1 _4584_/X sky130_fd_sc_hd__clkbuf_4
Xinput51 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__buf_4
Xinput62 wbs_data_i[17] vssd1 vssd1 vccd1 vccd1 _5012_/A sky130_fd_sc_hd__buf_4
Xinput73 wbs_data_i[27] vssd1 vssd1 vccd1 vccd1 _5035_/A sky130_fd_sc_hd__buf_4
X_7372_ _7372_/CLK _7372_/D vssd1 vssd1 vccd1 vccd1 _7372_/Q sky130_fd_sc_hd__dfxtp_1
X_3535_ _3534_/X _7710_/Q _3535_/S vssd1 vssd1 vccd1 vccd1 _3536_/A sky130_fd_sc_hd__mux2_1
Xinput84 wbs_data_i[8] vssd1 vssd1 vccd1 vccd1 _4993_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6254_ _6254_/A vssd1 vssd1 vccd1 vccd1 _6254_/X sky130_fd_sc_hd__buf_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5205_ _5205_/A vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5136_ _7130_/Q _7053_/Q _7045_/Q _7266_/Q _5132_/X _5135_/X vssd1 vssd1 vccd1 vccd1
+ _5136_/X sky130_fd_sc_hd__mux4_1
X_5067_ _5067_/A vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__clkbuf_1
X_4018_ _4018_/A vssd1 vssd1 vccd1 vccd1 _7489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5969_ _5901_/S _5962_/Y _5964_/Y _5966_/Y _5968_/Y vssd1 vssd1 vccd1 vccd1 _5969_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7708_ _7708_/CLK _7708_/D vssd1 vssd1 vccd1 vccd1 _7708_/Q sky130_fd_sc_hd__dfxtp_1
X_7639_ _7731_/CLK _7639_/D vssd1 vssd1 vccd1 vccd1 _7639_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2718_ _5707_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2718_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__3112_ clkbuf_0__3112_/X vssd1 vssd1 vccd1 vccd1 _6618__74/A sky130_fd_sc_hd__clkbuf_16
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6872_ _6870_/X _6872_/B _6872_/C vssd1 vssd1 vccd1 vccd1 _6873_/A sky130_fd_sc_hd__and3b_1
X_5823_ _5856_/A vssd1 vssd1 vccd1 vccd1 _5823_/X sky130_fd_sc_hd__buf_4
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5754_ _4997_/A _7188_/Q _5758_/S vssd1 vssd1 vccd1 vccd1 _5755_/A sky130_fd_sc_hd__mux2_1
X_4705_ _4705_/A vssd1 vssd1 vccd1 vccd1 _7182_/D sky130_fd_sc_hd__clkbuf_1
X_4636_ _4255_/X _7244_/Q _4640_/S vssd1 vssd1 vccd1 vccd1 _4637_/A sky130_fd_sc_hd__mux2_1
X_7424_ _7424_/CLK _7424_/D vssd1 vssd1 vccd1 vccd1 _7424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7355_ _7355_/CLK _7355_/D vssd1 vssd1 vccd1 vccd1 _7355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4567_ _4566_/X _7272_/Q _4576_/S vssd1 vssd1 vccd1 vccd1 _4568_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3518_ _3547_/S vssd1 vssd1 vccd1 vccd1 _3535_/S sky130_fd_sc_hd__clkbuf_2
X_7286_ _7286_/CLK _7286_/D vssd1 vssd1 vccd1 vccd1 _7286_/Q sky130_fd_sc_hd__dfxtp_1
X_4498_ _4226_/X _7305_/Q _4498_/S vssd1 vssd1 vccd1 vccd1 _4499_/A sky130_fd_sc_hd__mux2_1
X_6237_ _6237_/A vssd1 vssd1 vccd1 vccd1 _7330_/D sky130_fd_sc_hd__clkbuf_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6803_/B _6781_/A vssd1 vssd1 vccd1 vccd1 _6768_/A sky130_fd_sc_hd__or2_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _7081_/Q _7082_/Q _5585_/B _5185_/B vssd1 vssd1 vccd1 vccd1 _5380_/B sky130_fd_sc_hd__o31a_2
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6099_ _6450_/B _6139_/B _6093_/Y _6098_/Y vssd1 vssd1 vccd1 vccd1 _6492_/C sky130_fd_sc_hd__a31o_1
XFILLER_72_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6178__360 _6180__362/A vssd1 vssd1 vccd1 vccd1 _7290_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6042__324 _6042__324/A vssd1 vssd1 vccd1 vccd1 _7250_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5470_ _5458_/X _7194_/Q input10/X _5102_/D vssd1 vssd1 vccd1 vccd1 _5470_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4421_ _4421_/A vssd1 vssd1 vccd1 vccd1 _7338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7140_ _7140_/CLK _7140_/D vssd1 vssd1 vccd1 vccd1 _7140_/Q sky130_fd_sc_hd__dfxtp_1
X_4352_ _4782_/S vssd1 vssd1 vccd1 vccd1 _4774_/S sky130_fd_sc_hd__clkbuf_4
X_4283_ _4283_/A _4642_/A vssd1 vssd1 vccd1 vccd1 _4299_/S sky130_fd_sc_hd__or2_1
X_7071_ _7516_/CLK _7071_/D vssd1 vssd1 vccd1 vccd1 _7071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924_ _6924_/A vssd1 vssd1 vccd1 vccd1 _7674_/D sky130_fd_sc_hd__clkbuf_1
X_6855_ _6868_/A _6855_/B _6855_/C vssd1 vssd1 vccd1 vccd1 _6856_/A sky130_fd_sc_hd__and3_1
X_3998_ _3664_/X _7518_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _3999_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6786_ _5281_/X _6816_/A _6098_/Y _7650_/Q vssd1 vssd1 vccd1 vccd1 _6788_/B sky130_fd_sc_hd__o2bb2a_1
X_5737_ _6260_/A vssd1 vssd1 vccd1 vccd1 _5737_/X sky130_fd_sc_hd__buf_1
XFILLER_108_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7407_ _7407_/CLK _7407_/D vssd1 vssd1 vccd1 vccd1 _7407_/Q sky130_fd_sc_hd__dfxtp_1
X_4619_ _4619_/A vssd1 vssd1 vccd1 vccd1 _7252_/D sky130_fd_sc_hd__clkbuf_1
X_5599_ _5599_/A vssd1 vssd1 vccd1 vccd1 _7083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7338_ _7338_/CLK _7338_/D vssd1 vssd1 vccd1 vccd1 _7338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7269_ _7269_/CLK _7269_/D vssd1 vssd1 vccd1 vccd1 _7269_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_31 _5049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_20 _7308_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_42 _6919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_86 _3813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_53 _3801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_75 _7437_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_64 _5482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3094_ clkbuf_0__3094_/X vssd1 vssd1 vccd1 vccd1 _6356__484/A sky130_fd_sc_hd__clkbuf_16
XFILLER_119_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4970_ _5766_/A _4979_/B vssd1 vssd1 vccd1 vccd1 _4971_/A sky130_fd_sc_hd__and2_1
X_3921_ _3920_/X _7551_/Q _3924_/S vssd1 vssd1 vccd1 vccd1 _3922_/A sky130_fd_sc_hd__mux2_1
X_3852_ _3744_/X _7577_/Q _3852_/S vssd1 vssd1 vccd1 vccd1 _3853_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6571_ _6571_/A _6571_/B vssd1 vssd1 vccd1 vccd1 _6577_/B sky130_fd_sc_hd__nor2_1
X_3783_ _3783_/A vssd1 vssd1 vccd1 vccd1 _7603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5453_ _7722_/Q vssd1 vssd1 vccd1 vccd1 _6129_/A sky130_fd_sc_hd__buf_4
X_5384_ _7705_/Q _4396_/X _5383_/X vssd1 vssd1 vccd1 vccd1 _5384_/X sky130_fd_sc_hd__o21a_1
X_4404_ _7345_/Q _4325_/X _4410_/S vssd1 vssd1 vccd1 vccd1 _4405_/A sky130_fd_sc_hd__mux2_1
XCaravelHost_198 vssd1 vssd1 vccd1 vccd1 CaravelHost_198/HI core0Index[5] sky130_fd_sc_hd__conb_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7123_ _7123_/CLK _7123_/D vssd1 vssd1 vccd1 vccd1 _7123_/Q sky130_fd_sc_hd__dfxtp_1
X_4335_ _7363_/Q _4334_/X _4335_/S vssd1 vssd1 vccd1 vccd1 _4336_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7054_ _7054_/CLK _7054_/D vssd1 vssd1 vccd1 vccd1 _7054_/Q sky130_fd_sc_hd__dfxtp_1
X_4266_ _4281_/S vssd1 vssd1 vccd1 vccd1 _4275_/S sky130_fd_sc_hd__clkbuf_2
X_6005_ _6005_/A _6005_/B vssd1 vssd1 vccd1 vccd1 _6005_/Y sky130_fd_sc_hd__nor2_1
X_4197_ _4100_/X _7414_/Q _4203_/S vssd1 vssd1 vccd1 vccd1 _4198_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2966_ _6080_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2966_/X sky130_fd_sc_hd__clkbuf_16
X_6907_ _6921_/C vssd1 vssd1 vccd1 vccd1 _6923_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6430__62 _6432__64/A vssd1 vssd1 vccd1 vccd1 _7484_/CLK sky130_fd_sc_hd__inv_2
X_6838_ _7647_/Q vssd1 vssd1 vccd1 vccd1 _6847_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6769_ _7658_/Q vssd1 vssd1 vccd1 vccd1 _6878_/A sky130_fd_sc_hd__inv_2
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6949__38 _6950__39/A vssd1 vssd1 vccd1 vccd1 _7694_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3291_ clkbuf_0__3291_/X vssd1 vssd1 vccd1 vccd1 _6932_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3077_ clkbuf_0__3077_/X vssd1 vssd1 vccd1 vccd1 _6264__411/A sky130_fd_sc_hd__clkbuf_16
XFILLER_69_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4120_ _4120_/A vssd1 vssd1 vccd1 vccd1 _7448_/D sky130_fd_sc_hd__clkbuf_1
X_4051_ _4051_/A vssd1 vssd1 vccd1 vccd1 _7475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 caravel_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_4
XFILLER_110_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4953_ _4953_/A vssd1 vssd1 vccd1 vccd1 _7036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3904_ _3904_/A vssd1 vssd1 vccd1 vccd1 _7557_/D sky130_fd_sc_hd__clkbuf_1
X_7672_ _7674_/CLK _7672_/D vssd1 vssd1 vccd1 vccd1 _7672_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4884_ _4820_/X _7079_/Q _4892_/S vssd1 vssd1 vccd1 vccd1 _4885_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3835_ _3835_/A vssd1 vssd1 vccd1 vccd1 _7585_/D sky130_fd_sc_hd__clkbuf_1
X_3766_ _3652_/X _7610_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3767_/A sky130_fd_sc_hd__mux2_1
X_6554_ _6553_/B _6553_/C _6558_/B vssd1 vssd1 vccd1 vccd1 _6555_/C sky130_fd_sc_hd__a21o_1
X_5505_ _5706_/A vssd1 vssd1 vccd1 vccd1 _5505_/X sky130_fd_sc_hd__buf_1
X_6485_ _6486_/B _6486_/C _6541_/B vssd1 vssd1 vccd1 vccd1 _6485_/X sky130_fd_sc_hd__a21bo_1
X_3697_ _3526_/X _7635_/Q _3701_/S vssd1 vssd1 vccd1 vccd1 _3698_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5436_ _5494_/S _5436_/B _5436_/C vssd1 vssd1 vccd1 vccd1 _5436_/X sky130_fd_sc_hd__and3_1
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5367_ _5349_/S _5366_/X _5178_/A vssd1 vssd1 vccd1 vccd1 _5367_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5298_ _7545_/Q _7435_/Q _7403_/Q _7387_/Q _4381_/A _5252_/X vssd1 vssd1 vccd1 vccd1
+ _5298_/X sky130_fd_sc_hd__mux4_1
X_7106_ _7106_/CLK _7106_/D vssd1 vssd1 vccd1 vccd1 _7106_/Q sky130_fd_sc_hd__dfxtp_1
X_5697__252 _5699__254/A vssd1 vssd1 vccd1 vccd1 _7146_/CLK sky130_fd_sc_hd__inv_2
X_4318_ _4235_/X _7368_/Q _4318_/S vssd1 vssd1 vccd1 vccd1 _4319_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7037_ _7037_/CLK _7037_/D vssd1 vssd1 vccd1 vccd1 _7037_/Q sky130_fd_sc_hd__dfxtp_1
X_4249_ _7671_/Q vssd1 vssd1 vccd1 vccd1 _4249_/X sky130_fd_sc_hd__buf_2
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3096_ _6358_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3096_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2715_ clkbuf_0__2715_/X vssd1 vssd1 vccd1 vccd1 _5699__254/A sky130_fd_sc_hd__clkbuf_16
XFILLER_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3620_ _3526_/X _7696_/Q _3624_/S vssd1 vssd1 vccd1 vccd1 _3621_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__3274_ clkbuf_0__3274_/X vssd1 vssd1 vccd1 vccd1 _6662__108/A sky130_fd_sc_hd__clkbuf_16
X_3551_ _3983_/B vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3482_ _3484_/A _3484_/B _3481_/X vssd1 vssd1 vccd1 vccd1 _3483_/B sky130_fd_sc_hd__a21oi_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5221_ _5257_/A _5220_/X _5178_/X vssd1 vssd1 vccd1 vccd1 _5221_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5152_ _5213_/A vssd1 vssd1 vccd1 vccd1 _5163_/A sky130_fd_sc_hd__clkbuf_2
X_4103_ _7672_/Q vssd1 vssd1 vccd1 vccd1 _4103_/X sky130_fd_sc_hd__clkbuf_2
X_5083_ _5083_/A vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4034_ _4034_/A vssd1 vssd1 vccd1 vccd1 _7482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5985_ _6005_/A _5985_/B vssd1 vssd1 vccd1 vccd1 _5985_/Y sky130_fd_sc_hd__nor2_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7724_ _7731_/CLK _7724_/D vssd1 vssd1 vccd1 vccd1 _7724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4936_ _4936_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4952_/S sky130_fd_sc_hd__nand2_1
X_7655_ _7655_/CLK _7655_/D vssd1 vssd1 vccd1 vccd1 _7655_/Q sky130_fd_sc_hd__dfxtp_1
X_4867_ _4867_/A vssd1 vssd1 vccd1 vccd1 _7113_/D sky130_fd_sc_hd__clkbuf_1
X_3818_ _3818_/A vssd1 vssd1 vccd1 vccd1 _7591_/D sky130_fd_sc_hd__clkbuf_1
X_7586_ _7586_/CLK _7586_/D vssd1 vssd1 vccd1 vccd1 _7586_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2665_ _5579_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2665_/X sky130_fd_sc_hd__clkbuf_16
X_6606_ _6556_/B _6567_/A _6604_/Y _6464_/Y vssd1 vssd1 vccd1 vccd1 _6606_/X sky130_fd_sc_hd__a211o_1
X_4798_ _7139_/Q _4581_/A _4800_/S vssd1 vssd1 vccd1 vccd1 _4799_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6537_ _6567_/A vssd1 vssd1 vccd1 vccd1 _6562_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3749_ _3749_/A vssd1 vssd1 vccd1 vccd1 _7616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6468_ _7506_/Q vssd1 vssd1 vccd1 vccd1 _6571_/A sky130_fd_sc_hd__inv_2
Xoutput150 _4989_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[6] sky130_fd_sc_hd__buf_2
Xoutput161 _5195_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[0] sky130_fd_sc_hd__buf_2
X_5419_ _5413_/A _5416_/X _5418_/X _4368_/A vssd1 vssd1 vccd1 vccd1 _5419_/X sky130_fd_sc_hd__o211a_1
XFILLER_114_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput183 _5279_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput172 _5240_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[1] sky130_fd_sc_hd__buf_2
XFILLER_101_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2629_ clkbuf_0__2629_/X vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5770_ _5012_/A _7195_/Q _5776_/S vssd1 vssd1 vccd1 vccd1 _5771_/A sky130_fd_sc_hd__mux2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4721_/A vssd1 vssd1 vccd1 vccd1 _7175_/D sky130_fd_sc_hd__clkbuf_1
X_4652_ _4252_/X _7237_/Q _4652_/S vssd1 vssd1 vccd1 vccd1 _4653_/A sky130_fd_sc_hd__mux2_1
X_7440_ _7440_/CLK _7440_/D vssd1 vssd1 vccd1 vccd1 _7440_/Q sky130_fd_sc_hd__dfxtp_1
Xinput30 caravel_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_4
X_3603_ _7321_/Q vssd1 vssd1 vccd1 vccd1 _3603_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4583_ _4583_/A vssd1 vssd1 vccd1 vccd1 _7267_/D sky130_fd_sc_hd__clkbuf_1
Xinput41 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__buf_4
Xinput63 wbs_data_i[18] vssd1 vssd1 vccd1 vccd1 _5016_/A sky130_fd_sc_hd__buf_4
Xinput52 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__buf_4
X_7371_ _7371_/CLK _7371_/D vssd1 vssd1 vccd1 vccd1 _7371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3534_ _3914_/A vssd1 vssd1 vccd1 vccd1 _3534_/X sky130_fd_sc_hd__buf_2
Xinput85 wbs_data_i[9] vssd1 vssd1 vccd1 vccd1 _4995_/A sky130_fd_sc_hd__buf_4
Xinput74 wbs_data_i[28] vssd1 vssd1 vccd1 vccd1 _5038_/A sky130_fd_sc_hd__buf_4
Xclkbuf_4_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7670_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_103_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5204_ _7527_/Q _7107_/Q _7559_/Q _7123_/Q _5132_/X _5135_/X vssd1 vssd1 vccd1 vccd1
+ _5204_/X sky130_fd_sc_hd__mux4_1
X_6746__176 _6747__177/A vssd1 vssd1 vccd1 vccd1 _7620_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5135_ _5285_/S vssd1 vssd1 vccd1 vccd1 _5135_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5066_ _5066_/A _5068_/B vssd1 vssd1 vccd1 vccd1 _5067_/A sky130_fd_sc_hd__and2_1
X_4017_ _7489_/Q _3600_/X _4019_/S vssd1 vssd1 vccd1 vccd1 _4018_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5968_ _5923_/A _5967_/X _5929_/X vssd1 vssd1 vccd1 vccd1 _5968_/Y sky130_fd_sc_hd__o21ai_1
X_6621__76 _6621__76/A vssd1 vssd1 vccd1 vccd1 _7519_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7707_ _7707_/CLK _7707_/D vssd1 vssd1 vccd1 vccd1 _7707_/Q sky130_fd_sc_hd__dfxtp_1
X_4919_ _4934_/S vssd1 vssd1 vccd1 vccd1 _4928_/S sky130_fd_sc_hd__buf_2
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5899_ _5897_/X _5898_/X _5899_/S vssd1 vssd1 vccd1 vccd1 _5899_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_0__2717_ _5706_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2717_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7638_ _7731_/CLK _7638_/D vssd1 vssd1 vccd1 vccd1 _7638_/Q sky130_fd_sc_hd__dfxtp_1
X_7569_ _7569_/CLK _7569_/D vssd1 vssd1 vccd1 vccd1 _7569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__3111_ clkbuf_0__3111_/X vssd1 vssd1 vccd1 vccd1 _6438__69/A sky130_fd_sc_hd__clkbuf_16
XFILLER_112_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6871_ _7653_/Q _6870_/C _7654_/Q vssd1 vssd1 vccd1 vccd1 _6872_/C sky130_fd_sc_hd__a21o_1
Xclkbuf_1_0__f__2757_ clkbuf_0__2757_/X vssd1 vssd1 vccd1 vccd1 _5808__297/A sky130_fd_sc_hd__clkbuf_16
X_5822_ _7311_/Q vssd1 vssd1 vccd1 vccd1 _5908_/A sky130_fd_sc_hd__buf_4
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5753_ _5753_/A vssd1 vssd1 vccd1 vccd1 _7187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4704_ _4572_/X _7182_/Q _4706_/S vssd1 vssd1 vccd1 vccd1 _4705_/A sky130_fd_sc_hd__mux2_1
X_4635_ _4635_/A vssd1 vssd1 vccd1 vccd1 _7245_/D sky130_fd_sc_hd__clkbuf_1
X_7423_ _7423_/CLK _7423_/D vssd1 vssd1 vccd1 vccd1 _7423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4566_ _4566_/A vssd1 vssd1 vccd1 vccd1 _4566_/X sky130_fd_sc_hd__buf_2
X_7354_ _7354_/CLK _7354_/D vssd1 vssd1 vccd1 vccd1 _7354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3517_ _4283_/A _4121_/A vssd1 vssd1 vccd1 vccd1 _3547_/S sky130_fd_sc_hd__or2_2
XFILLER_103_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4497_ _4497_/A vssd1 vssd1 vccd1 vccd1 _7306_/D sky130_fd_sc_hd__clkbuf_1
X_7285_ _7731_/CLK _7285_/D vssd1 vssd1 vccd1 vccd1 _7285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6236_ _7525_/Q _6236_/B _6236_/C _7715_/Q vssd1 vssd1 vccd1 vccd1 _6237_/A sky130_fd_sc_hd__and4b_1
XFILLER_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _7638_/Q vssd1 vssd1 vccd1 vccd1 _6781_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5118_/A _5118_/B _5118_/C vssd1 vssd1 vccd1 vccd1 _5187_/A sky130_fd_sc_hd__or3_2
X_6437__68 _6437__68/A vssd1 vssd1 vccd1 vccd1 _7490_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6098_ _7721_/Q vssd1 vssd1 vccd1 vccd1 _6098_/Y sky130_fd_sc_hd__inv_2
X_5049_ _5049_/A _5057_/B vssd1 vssd1 vccd1 vccd1 _5050_/A sky130_fd_sc_hd__and2_1
XFILLER_85_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6371__495 _6375__499/A vssd1 vssd1 vccd1 vccd1 _7437_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4420_ _4211_/X _7338_/Q _4428_/S vssd1 vssd1 vccd1 vccd1 _4421_/A sky130_fd_sc_hd__mux2_1
X_4351_ _4562_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _4782_/S sky130_fd_sc_hd__nor2_2
XFILLER_98_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4282_ _4282_/A vssd1 vssd1 vccd1 vccd1 _7384_/D sky130_fd_sc_hd__clkbuf_1
X_7070_ _7190_/CLK _7070_/D vssd1 vssd1 vccd1 vccd1 _7070_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5691__247 _5691__247/A vssd1 vssd1 vccd1 vccd1 _7141_/CLK sky130_fd_sc_hd__inv_2
X_6923_ _6923_/A _6923_/B vssd1 vssd1 vccd1 vccd1 _6924_/A sky130_fd_sc_hd__and2_1
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6854_ _6863_/C _6857_/C vssd1 vssd1 vccd1 vccd1 _6855_/C sky130_fd_sc_hd__or2_1
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5805_ _6018_/A vssd1 vssd1 vccd1 vccd1 _5805_/X sky130_fd_sc_hd__buf_1
X_3997_ _3997_/A vssd1 vssd1 vccd1 vccd1 _7519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6785_ _6783_/Y _6784_/X _7655_/Q _6143_/A vssd1 vssd1 vccd1 vccd1 _6789_/B sky130_fd_sc_hd__a211o_1
X_4618_ _7252_/Q _3917_/A _4622_/S vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__mux2_1
X_7406_ _7406_/CLK _7406_/D vssd1 vssd1 vccd1 vccd1 _7406_/Q sky130_fd_sc_hd__dfxtp_2
X_5598_ _7083_/Q _5055_/A _5602_/S vssd1 vssd1 vccd1 vccd1 _5599_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6019__305 _6021__307/A vssd1 vssd1 vccd1 vccd1 _7231_/CLK sky130_fd_sc_hd__inv_2
X_4549_ _4549_/A vssd1 vssd1 vccd1 vccd1 _7282_/D sky130_fd_sc_hd__clkbuf_1
X_7337_ _7337_/CLK _7337_/D vssd1 vssd1 vccd1 vccd1 _7337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7268_ _7268_/CLK _7268_/D vssd1 vssd1 vccd1 vccd1 _7268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6219_ _6219_/A vssd1 vssd1 vccd1 vccd1 _7322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_10 _4328_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7199_ _7674_/CLK _7199_/D vssd1 vssd1 vccd1 vccd1 _7199_/Q sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_32 _5049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_43 _6919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_21 _7406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_54 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_65 _6119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_76 _7338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_87 _3819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3093_ clkbuf_0__3093_/X vssd1 vssd1 vccd1 vccd1 _6350__479/A sky130_fd_sc_hd__clkbuf_16
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6703__141 _6706__144/A vssd1 vssd1 vccd1 vccd1 _7585_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3920_ _3920_/A vssd1 vssd1 vccd1 vccd1 _3920_/X sky130_fd_sc_hd__buf_4
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3851_ _3851_/A vssd1 vssd1 vccd1 vccd1 _7578_/D sky130_fd_sc_hd__clkbuf_1
X_3782_ _3738_/X _7603_/Q _3786_/S vssd1 vssd1 vccd1 vccd1 _3783_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6570_ _6566_/X _6568_/X _6569_/X vssd1 vssd1 vccd1 vccd1 _7505_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5452_ _6137_/A _5448_/X _5449_/X _5451_/X vssd1 vssd1 vccd1 vccd1 _5452_/X sky130_fd_sc_hd__a31o_1
X_5383_ _5325_/S _7292_/Q _5148_/A vssd1 vssd1 vccd1 vccd1 _5383_/X sky130_fd_sc_hd__o21ba_1
X_4403_ _4403_/A vssd1 vssd1 vccd1 vccd1 _7346_/D sky130_fd_sc_hd__clkbuf_1
X_7122_ _7122_/CLK _7122_/D vssd1 vssd1 vccd1 vccd1 _7122_/Q sky130_fd_sc_hd__dfxtp_1
XCaravelHost_199 vssd1 vssd1 vccd1 vccd1 CaravelHost_199/HI core0Index[6] sky130_fd_sc_hd__conb_1
X_4334_ _7324_/Q vssd1 vssd1 vccd1 vccd1 _4334_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7053_ _7053_/CLK _7053_/D vssd1 vssd1 vccd1 vccd1 _7053_/Q sky130_fd_sc_hd__dfxtp_1
X_6004_ _7629_/Q _7621_/Q _7605_/Q _7597_/Q _5823_/X _5925_/X vssd1 vssd1 vccd1 vccd1
+ _6005_/B sky130_fd_sc_hd__mux4_2
XFILLER_86_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4265_ _4562_/A _4265_/B vssd1 vssd1 vccd1 vccd1 _4281_/S sky130_fd_sc_hd__nor2_2
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4196_ _4196_/A vssd1 vssd1 vccd1 vccd1 _7415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6906_ input1/X _6892_/X _6905_/X _6886_/X vssd1 vssd1 vccd1 vccd1 _7666_/D sky130_fd_sc_hd__o211a_1
X_6837_ _6837_/A vssd1 vssd1 vccd1 vccd1 _7646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6322__456 _6323__457/A vssd1 vssd1 vccd1 vccd1 _7398_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6768_ _6768_/A vssd1 vssd1 vccd1 vccd1 _6889_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5719_ _5725_/A vssd1 vssd1 vccd1 vccd1 _5719_/X sky130_fd_sc_hd__buf_1
XFILLER_108_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__3290_ clkbuf_0__3290_/X vssd1 vssd1 vccd1 vccd1 _6747__177/A sky130_fd_sc_hd__clkbuf_16
XFILLER_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3076_ clkbuf_0__3076_/X vssd1 vssd1 vccd1 vccd1 _6289_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4050_ _3914_/X _7475_/Q _4050_/S vssd1 vssd1 vccd1 vccd1 _4051_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 caravel_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4952_ _3819_/X _7036_/Q _4952_/S vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__mux2_1
X_3903_ _3899_/X _7557_/Q _3915_/S vssd1 vssd1 vccd1 vccd1 _3904_/A sky130_fd_sc_hd__mux2_1
X_7671_ _7674_/CLK _7671_/D vssd1 vssd1 vccd1 vccd1 _7671_/Q sky130_fd_sc_hd__dfxtp_2
X_4883_ _4898_/S vssd1 vssd1 vccd1 vccd1 _4892_/S sky130_fd_sc_hd__clkbuf_4
X_3834_ _3744_/X _7585_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3835_/A sky130_fd_sc_hd__mux2_1
X_3765_ _3765_/A vssd1 vssd1 vccd1 vccd1 _7611_/D sky130_fd_sc_hd__clkbuf_1
X_6553_ _6558_/B _6553_/B _6553_/C vssd1 vssd1 vccd1 vccd1 _6559_/B sky130_fd_sc_hd__and3_1
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3696_ _3696_/A vssd1 vssd1 vccd1 vccd1 _7636_/D sky130_fd_sc_hd__clkbuf_1
X_6484_ _7500_/Q vssd1 vssd1 vccd1 vccd1 _6541_/B sky130_fd_sc_hd__clkbuf_2
X_5435_ _5381_/Y _5420_/X _5433_/X _5441_/D _6476_/A vssd1 vssd1 vccd1 vccd1 _5436_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_99_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5366_ _7175_/Q _7307_/Q _7493_/Q _7183_/Q _5207_/A _5325_/S vssd1 vssd1 vccd1 vccd1
+ _5366_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4317_ _4317_/A vssd1 vssd1 vccd1 vccd1 _7369_/D sky130_fd_sc_hd__clkbuf_1
X_7105_ _7190_/CLK _7105_/D vssd1 vssd1 vccd1 vccd1 _7105_/Q sky130_fd_sc_hd__dfxtp_1
X_5297_ _5158_/X _5287_/X _5289_/Y _5296_/X _5161_/X vssd1 vssd1 vccd1 vccd1 _5308_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7036_ _7036_/CLK _7036_/D vssd1 vssd1 vccd1 vccd1 _7036_/Q sky130_fd_sc_hd__dfxtp_1
X_4248_ _4248_/A vssd1 vssd1 vccd1 vccd1 _7397_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3095_ _6357_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3095_/X sky130_fd_sc_hd__clkbuf_16
X_4179_ _4100_/X _7422_/Q _4185_/S vssd1 vssd1 vccd1 vccd1 _4180_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6954__42 _6955__43/A vssd1 vssd1 vccd1 vccd1 _7698_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6246__398 _6246__398/A vssd1 vssd1 vccd1 vccd1 _7338_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2714_ clkbuf_0__2714_/X vssd1 vssd1 vccd1 vccd1 _5691__247/A sky130_fd_sc_hd__clkbuf_16
XFILLER_19_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__3273_ clkbuf_0__3273_/X vssd1 vssd1 vccd1 vccd1 _6682_/A sky130_fd_sc_hd__clkbuf_16
X_3550_ _7356_/Q vssd1 vssd1 vccd1 vccd1 _3983_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_1__f__3059_ clkbuf_0__3059_/X vssd1 vssd1 vccd1 vccd1 _6240__393/A sky130_fd_sc_hd__clkbuf_16
X_3481_ _7318_/Q _5929_/A vssd1 vssd1 vccd1 vccd1 _3481_/X sky130_fd_sc_hd__xor2_1
X_5220_ _7369_/Q _7340_/Q _7332_/Q _7295_/Q _5138_/X _5293_/A vssd1 vssd1 vccd1 vccd1
+ _5220_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5151_ _7349_/Q vssd1 vssd1 vccd1 vccd1 _5213_/A sky130_fd_sc_hd__clkinv_2
X_5082_ _7194_/Q _5090_/B vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__and2_1
XFILLER_96_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4102_ _4102_/A vssd1 vssd1 vccd1 vccd1 _7454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4033_ _3917_/X _7482_/Q _4037_/S vssd1 vssd1 vccd1 vccd1 _4034_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5984_ _7628_/Q _7620_/Q _7604_/Q _7596_/Q _5823_/X _5925_/X vssd1 vssd1 vccd1 vccd1
+ _5985_/B sky130_fd_sc_hd__mux4_2
X_7723_ _7723_/CLK _7723_/D vssd1 vssd1 vccd1 vccd1 _7723_/Q sky130_fd_sc_hd__dfxtp_1
X_4935_ _4935_/A vssd1 vssd1 vccd1 vccd1 _7045_/D sky130_fd_sc_hd__clkbuf_1
X_7654_ _7655_/CLK _7654_/D vssd1 vssd1 vccd1 vccd1 _7654_/Q sky130_fd_sc_hd__dfxtp_1
X_4866_ _4820_/X _7113_/Q _4874_/S vssd1 vssd1 vccd1 vccd1 _4867_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3817_ _7591_/Q _3816_/X _3820_/S vssd1 vssd1 vccd1 vccd1 _3818_/A sky130_fd_sc_hd__mux2_1
X_7585_ _7585_/CLK _7585_/D vssd1 vssd1 vccd1 vccd1 _7585_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2664_ _5573_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2664_/X sky130_fd_sc_hd__clkbuf_16
X_4797_ _4797_/A vssd1 vssd1 vccd1 vccd1 _7140_/D sky130_fd_sc_hd__clkbuf_1
X_6605_ _6579_/B _6579_/C _6604_/Y vssd1 vssd1 vccd1 vccd1 _6605_/Y sky130_fd_sc_hd__a21oi_1
X_3748_ _3747_/X _7616_/Q _3754_/S vssd1 vssd1 vccd1 vccd1 _3749_/A sky130_fd_sc_hd__mux2_1
X_6536_ _6561_/A vssd1 vssd1 vccd1 vccd1 _6556_/B sky130_fd_sc_hd__clkbuf_2
X_3679_ _3679_/A vssd1 vssd1 vccd1 vccd1 _7680_/D sky130_fd_sc_hd__clkbuf_1
X_6467_ _6452_/A _6446_/B _6137_/A vssd1 vssd1 vccd1 vccd1 _6470_/C sky130_fd_sc_hd__o21ai_1
Xoutput140 _5034_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[26] sky130_fd_sc_hd__buf_2
Xoutput151 _4991_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[7] sky130_fd_sc_hd__buf_2
X_5418_ _5418_/A _5418_/B vssd1 vssd1 vccd1 vccd1 _5418_/X sky130_fd_sc_hd__or2_1
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6172__356 _6173__357/A vssd1 vssd1 vccd1 vccd1 _7286_/CLK sky130_fd_sc_hd__inv_2
X_5349_ _5347_/X _5348_/X _5349_/S vssd1 vssd1 vccd1 vccd1 _5349_/X sky130_fd_sc_hd__mux2_1
Xoutput162 _5455_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput173 _5478_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[20] sky130_fd_sc_hd__buf_2
Xoutput184 _5490_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7019_ _7003_/X _7019_/B vssd1 vssd1 vccd1 vccd1 _7020_/A sky130_fd_sc_hd__and2b_1
Xclkbuf_0__3078_ _6268_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3078_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6927__20 _6931__24/A vssd1 vssd1 vccd1 vccd1 _7676_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5712__264 _5712__264/A vssd1 vssd1 vccd1 vccd1 _7158_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6335__466 _6337__468/A vssd1 vssd1 vccd1 vccd1 _7408_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2628_ clkbuf_0__2628_/X vssd1 vssd1 vccd1 vccd1 _5502__182/A sky130_fd_sc_hd__clkbuf_16
X_6659__105 _6662__108/A vssd1 vssd1 vccd1 vccd1 _7549_/CLK sky130_fd_sc_hd__inv_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4569_/X _7175_/Q _4724_/S vssd1 vssd1 vccd1 vccd1 _4721_/A sky130_fd_sc_hd__mux2_1
X_4651_ _4651_/A vssd1 vssd1 vccd1 vccd1 _7238_/D sky130_fd_sc_hd__clkbuf_1
Xinput20 caravel_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_2
Xinput31 caravel_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
X_3602_ _3602_/A vssd1 vssd1 vccd1 vccd1 _7700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4582_ _4581_/X _7267_/Q _4585_/S vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__mux2_1
X_7370_ _7370_/CLK _7370_/D vssd1 vssd1 vccd1 vccd1 _7370_/Q sky130_fd_sc_hd__dfxtp_1
Xinput42 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__buf_4
Xinput53 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _5555_/B sky130_fd_sc_hd__buf_4
Xinput64 wbs_data_i[19] vssd1 vssd1 vccd1 vccd1 _5018_/A sky130_fd_sc_hd__buf_4
X_3533_ _7670_/Q vssd1 vssd1 vccd1 vccd1 _3914_/A sky130_fd_sc_hd__buf_2
Xinput86 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _5536_/A sky130_fd_sc_hd__buf_6
Xinput75 wbs_data_i[29] vssd1 vssd1 vccd1 vccd1 _5040_/A sky130_fd_sc_hd__buf_4
XFILLER_107_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6183_ _6195_/A vssd1 vssd1 vccd1 vccd1 _6183_/X sky130_fd_sc_hd__buf_1
X_5203_ _4375_/A _5202_/X _5163_/A vssd1 vssd1 vccd1 vccd1 _5203_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5134_ _5270_/A vssd1 vssd1 vccd1 vccd1 _5285_/S sky130_fd_sc_hd__clkbuf_4
X_5065_ _5065_/A vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__clkbuf_1
X_5655__218 _5655__218/A vssd1 vssd1 vccd1 vccd1 _7112_/CLK sky130_fd_sc_hd__inv_2
X_4016_ _4016_/A vssd1 vssd1 vccd1 vccd1 _7490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5967_ _7413_/Q _7381_/Q _7712_/Q _7635_/Q _5921_/X _5884_/X vssd1 vssd1 vccd1 vccd1
+ _5967_/X sky130_fd_sc_hd__mux4_1
X_7706_ _7706_/CLK _7706_/D vssd1 vssd1 vccd1 vccd1 _7706_/Q sky130_fd_sc_hd__dfxtp_1
X_4918_ _4918_/A _4918_/B vssd1 vssd1 vccd1 vccd1 _4934_/S sky130_fd_sc_hd__nor2_2
XFILLER_21_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5898_ _7244_/Q _7228_/Q _7474_/Q _7466_/Q _5908_/A _5823_/X vssd1 vssd1 vccd1 vccd1
+ _5898_/X sky130_fd_sc_hd__mux4_1
X_7637_ _7637_/CLK _7637_/D vssd1 vssd1 vccd1 vccd1 _7637_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2716_ _5700_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2716_/X sky130_fd_sc_hd__clkbuf_16
X_4849_ _4849_/A vssd1 vssd1 vccd1 vccd1 _7121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7568_ _7568_/CLK _7568_/D vssd1 vssd1 vccd1 vccd1 _7568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7499_ _7652_/CLK _7499_/D vssd1 vssd1 vccd1 vccd1 _7499_/Q sky130_fd_sc_hd__dfxtp_1
X_6519_ _6519_/A vssd1 vssd1 vccd1 vccd1 _7496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__3110_ clkbuf_0__3110_/X vssd1 vssd1 vccd1 vccd1 _6429__61/A sky130_fd_sc_hd__clkbuf_16
XFILLER_8_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5574__205 _5576__207/A vssd1 vssd1 vccd1 vccd1 _7073_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6870_ _7654_/Q _7653_/Q _6870_/C vssd1 vssd1 vccd1 vccd1 _6870_/X sky130_fd_sc_hd__and3_1
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5821_ _5959_/S _5821_/B vssd1 vssd1 vccd1 vccd1 _5821_/X sky130_fd_sc_hd__or2_1
XFILLER_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5752_ _4995_/A _7187_/Q _5758_/S vssd1 vssd1 vccd1 vccd1 _5753_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4703_ _4703_/A vssd1 vssd1 vccd1 vccd1 _7183_/D sky130_fd_sc_hd__clkbuf_1
X_4634_ _4252_/X _7245_/Q _4634_/S vssd1 vssd1 vccd1 vccd1 _4635_/A sky130_fd_sc_hd__mux2_1
X_7422_ _7422_/CLK _7422_/D vssd1 vssd1 vccd1 vccd1 _7422_/Q sky130_fd_sc_hd__dfxtp_1
X_4565_ _4565_/A vssd1 vssd1 vccd1 vccd1 _7273_/D sky130_fd_sc_hd__clkbuf_1
X_7353_ _7353_/CLK _7353_/D vssd1 vssd1 vccd1 vccd1 _7353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3516_ _3671_/A _4436_/A _3711_/C vssd1 vssd1 vccd1 vccd1 _4121_/A sky130_fd_sc_hd__nand3_4
X_7284_ _7284_/CLK _7284_/D vssd1 vssd1 vccd1 vccd1 _7284_/Q sky130_fd_sc_hd__dfxtp_1
X_4496_ _4223_/X _7306_/Q _4498_/S vssd1 vssd1 vccd1 vccd1 _4497_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6235_ _6235_/A vssd1 vssd1 vccd1 vccd1 _7329_/D sky130_fd_sc_hd__clkbuf_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _7639_/Q vssd1 vssd1 vccd1 vccd1 _6803_/B sky130_fd_sc_hd__inv_2
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6149_/A _6133_/A _6476_/A _6481_/A vssd1 vssd1 vccd1 vccd1 _6139_/B sky130_fd_sc_hd__nor4_1
X_5117_ _7101_/Q _7102_/Q _7092_/Q _7091_/Q vssd1 vssd1 vccd1 vccd1 _5118_/C sky130_fd_sc_hd__or4b_1
X_5048_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5057_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_111_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5516__188 _5517__189/A vssd1 vssd1 vccd1 vccd1 _7045_/CLK sky130_fd_sc_hd__inv_2
X_6999_ _6999_/A vssd1 vssd1 vccd1 vccd1 _7721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2962_ clkbuf_0__2962_/X vssd1 vssd1 vccd1 vccd1 _6079__349/A sky130_fd_sc_hd__clkbuf_16
XFILLER_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6185__366 _6186__367/A vssd1 vssd1 vccd1 vccd1 _7296_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4350_ _4350_/A _4350_/B vssd1 vssd1 vccd1 vccd1 _4356_/B sky130_fd_sc_hd__nand2_1
X_4281_ _7384_/Q _3603_/X _4281_/S vssd1 vssd1 vccd1 vccd1 _4282_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6922_ _6922_/A vssd1 vssd1 vccd1 vccd1 _7673_/D sky130_fd_sc_hd__clkbuf_1
X_6442__72 _6618__74/A vssd1 vssd1 vccd1 vccd1 _7494_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6853_ _6863_/C _6857_/C vssd1 vssd1 vccd1 vccd1 _6855_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3996_ _3660_/X _7519_/Q _4000_/S vssd1 vssd1 vccd1 vccd1 _3997_/A sky130_fd_sc_hd__mux2_1
X_6784_ _6784_/A _7643_/Q vssd1 vssd1 vccd1 vccd1 _6784_/X sky130_fd_sc_hd__or2_1
XFILLER_13_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4617_ _4617_/A vssd1 vssd1 vccd1 vccd1 _7253_/D sky130_fd_sc_hd__clkbuf_1
X_7405_ _7405_/CLK _7405_/D vssd1 vssd1 vccd1 vccd1 _7405_/Q sky130_fd_sc_hd__dfxtp_2
X_5597_ _5597_/A vssd1 vssd1 vccd1 vccd1 _7082_/D sky130_fd_sc_hd__clkbuf_1
X_4548_ _7282_/Q _3908_/A _4552_/S vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__mux2_1
X_7336_ _7336_/CLK _7336_/D vssd1 vssd1 vccd1 vccd1 _7336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7267_ _7267_/CLK _7267_/D vssd1 vssd1 vccd1 vccd1 _7267_/Q sky130_fd_sc_hd__dfxtp_1
X_4479_ _4473_/B _4479_/B _4486_/C vssd1 vssd1 vccd1 vccd1 _4480_/A sky130_fd_sc_hd__and3b_1
X_6218_ _7660_/Q _6220_/B vssd1 vssd1 vccd1 vccd1 _6219_/A sky130_fd_sc_hd__and2_1
X_7198_ _7727_/CLK _7198_/D vssd1 vssd1 vccd1 vccd1 _7198_/Q sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_33 _5049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_22 _7406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6149_ _6149_/A _7726_/Q vssd1 vssd1 vccd1 vccd1 _6483_/C sky130_fd_sc_hd__nor2_2
XINSDIODE2_11 _4337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_55 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_77 _7073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_66 _6137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_44 _6919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_88 _4217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3092_ clkbuf_0__3092_/X vssd1 vssd1 vccd1 vccd1 _6342__472/A sky130_fd_sc_hd__clkbuf_16
XFILLER_70_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3850_ _3741_/X _7578_/Q _3852_/S vssd1 vssd1 vccd1 vccd1 _3851_/A sky130_fd_sc_hd__mux2_1
X_3781_ _3781_/A vssd1 vssd1 vccd1 vccd1 _7604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5451_ _5444_/X _7187_/Q _5450_/X input34/X vssd1 vssd1 vccd1 vccd1 _5451_/X sky130_fd_sc_hd__a22o_1
X_5382_ _7078_/Q _7366_/Q _5397_/S vssd1 vssd1 vccd1 vccd1 _5382_/X sky130_fd_sc_hd__mux2_1
X_4402_ _7346_/Q _4320_/X _4410_/S vssd1 vssd1 vccd1 vccd1 _4403_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7121_ _7121_/CLK _7121_/D vssd1 vssd1 vccd1 vccd1 _7121_/Q sky130_fd_sc_hd__dfxtp_1
X_4333_ _4333_/A vssd1 vssd1 vccd1 vccd1 _7364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7052_ _7052_/CLK _7052_/D vssd1 vssd1 vccd1 vccd1 _7052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4264_ _4821_/A vssd1 vssd1 vccd1 vccd1 _4562_/A sky130_fd_sc_hd__buf_4
X_6003_ _6003_/A _6003_/B vssd1 vssd1 vccd1 vccd1 _6003_/Y sky130_fd_sc_hd__nor2_1
X_4195_ _4094_/X _7415_/Q _4203_/S vssd1 vssd1 vccd1 vccd1 _4196_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6905_ _7666_/Q _6905_/B vssd1 vssd1 vccd1 vccd1 _6905_/X sky130_fd_sc_hd__or2_1
X_6836_ _6843_/C _6836_/B _6859_/C vssd1 vssd1 vccd1 vccd1 _6837_/A sky130_fd_sc_hd__and3b_1
XFILLER_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3979_ _3664_/X _7527_/Q _3981_/S vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7319_ _7319_/CLK _7319_/D vssd1 vssd1 vccd1 vccd1 _7319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3075_ clkbuf_0__3075_/X vssd1 vssd1 vccd1 vccd1 _6388_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput7 caravel_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4951_ _4951_/A vssd1 vssd1 vccd1 vccd1 _7037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3902_ _3924_/S vssd1 vssd1 vccd1 vccd1 _3915_/S sky130_fd_sc_hd__clkbuf_2
X_7670_ _7670_/CLK _7670_/D vssd1 vssd1 vccd1 vccd1 _7670_/Q sky130_fd_sc_hd__dfxtp_2
X_4882_ _4882_/A _4900_/A vssd1 vssd1 vccd1 vccd1 _4898_/S sky130_fd_sc_hd__or2_2
X_3833_ _3833_/A vssd1 vssd1 vccd1 vccd1 _7586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3764_ _3648_/X _7611_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3765_/A sky130_fd_sc_hd__mux2_1
X_6552_ _6550_/X _6551_/X _6539_/X vssd1 vssd1 vccd1 vccd1 _7502_/D sky130_fd_sc_hd__o21a_1
X_3695_ _3522_/X _7636_/Q _3701_/S vssd1 vssd1 vccd1 vccd1 _3696_/A sky130_fd_sc_hd__mux2_1
X_6483_ _6483_/A _6483_/B _6483_/C _6483_/D vssd1 vssd1 vccd1 vccd1 _6483_/Y sky130_fd_sc_hd__nand4_1
XFILLER_118_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5434_ _7725_/Q vssd1 vssd1 vccd1 vccd1 _6476_/A sky130_fd_sc_hd__buf_4
XFILLER_105_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7104_ _7732_/CLK _7104_/D vssd1 vssd1 vccd1 vccd1 _7104_/Q sky130_fd_sc_hd__dfxtp_1
X_5365_ _5365_/A _5364_/X vssd1 vssd1 vccd1 vccd1 _5365_/X sky130_fd_sc_hd__or2b_1
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4316_ _4232_/X _7369_/Q _4318_/S vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__mux2_1
X_5296_ _5356_/A _5291_/Y _5293_/X _5295_/Y vssd1 vssd1 vccd1 vccd1 _5296_/X sky130_fd_sc_hd__a31o_1
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4247_ _4246_/X _7397_/Q _4253_/S vssd1 vssd1 vccd1 vccd1 _4248_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3094_ _6351_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3094_/X sky130_fd_sc_hd__clkbuf_16
X_7035_ _7035_/A vssd1 vssd1 vccd1 vccd1 _7732_/D sky130_fd_sc_hd__clkbuf_1
X_4178_ _4178_/A vssd1 vssd1 vccd1 vccd1 _7423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6819_ _6821_/A _7642_/Q _7641_/Q _6819_/D vssd1 vssd1 vccd1 vccd1 _6833_/D sky130_fd_sc_hd__and4_1
X_6652__100 _6656__104/A vssd1 vssd1 vccd1 vccd1 _7544_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2713_ clkbuf_0__2713_/X vssd1 vssd1 vccd1 vccd1 _5686__243/A sky130_fd_sc_hd__clkbuf_16
XFILLER_76_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6264__411 _6264__411/A vssd1 vssd1 vccd1 vccd1 _7351_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__3272_ clkbuf_0__3272_/X vssd1 vssd1 vccd1 vccd1 _6656__104/A sky130_fd_sc_hd__clkbuf_16
X_3480_ _7313_/Q vssd1 vssd1 vccd1 vccd1 _5929_/A sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__3058_ clkbuf_0__3058_/X vssd1 vssd1 vccd1 vccd1 _6213__389/A sky130_fd_sc_hd__clkbuf_16
XFILLER_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5150_ _5289_/A _5150_/B vssd1 vssd1 vccd1 vccd1 _5150_/X sky130_fd_sc_hd__or2_1
X_5081_ _5092_/A vssd1 vssd1 vccd1 vccd1 _5090_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4101_ _4100_/X _7454_/Q _4110_/S vssd1 vssd1 vccd1 vccd1 _4102_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4032_ _4032_/A vssd1 vssd1 vccd1 vccd1 _7483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5983_ _6003_/A _5983_/B vssd1 vssd1 vccd1 vccd1 _5983_/Y sky130_fd_sc_hd__nor2_1
X_4934_ _7045_/Q _4584_/A _4934_/S vssd1 vssd1 vccd1 vccd1 _4935_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7722_ _7722_/CLK _7722_/D vssd1 vssd1 vccd1 vccd1 _7722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7653_ _7655_/CLK _7653_/D vssd1 vssd1 vccd1 vccd1 _7653_/Q sky130_fd_sc_hd__dfxtp_1
X_4865_ _4880_/S vssd1 vssd1 vccd1 vccd1 _4874_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_33_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7584_ _7584_/CLK _7584_/D vssd1 vssd1 vccd1 vccd1 _7584_/Q sky130_fd_sc_hd__dfxtp_1
X_3816_ _7668_/Q vssd1 vssd1 vccd1 vccd1 _3816_/X sky130_fd_sc_hd__buf_6
X_4796_ _7140_/Q _4578_/A _4800_/S vssd1 vssd1 vccd1 vccd1 _4797_/A sky130_fd_sc_hd__mux2_1
X_6604_ _7512_/Q _7511_/Q _6604_/C vssd1 vssd1 vccd1 vccd1 _6604_/Y sky130_fd_sc_hd__nand3_1
X_6716__152 _6716__152/A vssd1 vssd1 vccd1 vccd1 _7596_/CLK sky130_fd_sc_hd__inv_2
X_3747_ _3917_/A vssd1 vssd1 vccd1 vccd1 _3747_/X sky130_fd_sc_hd__buf_2
X_6535_ _6543_/B _6535_/B _6583_/C vssd1 vssd1 vccd1 vccd1 _6535_/X sky130_fd_sc_hd__and3b_1
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3678_ _3526_/X _7680_/Q _3682_/S vssd1 vssd1 vccd1 vccd1 _3679_/A sky130_fd_sc_hd__mux2_1
X_6466_ _6594_/A _6503_/B _6500_/A _6500_/B vssd1 vssd1 vccd1 vccd1 _6466_/Y sky130_fd_sc_hd__o211ai_1
Xoutput141 _5036_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput130 _5013_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[17] sky130_fd_sc_hd__buf_2
Xoutput152 _4994_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[8] sky130_fd_sc_hd__buf_2
X_5417_ _7375_/Q _7346_/Q _7338_/Q _7301_/Q _5270_/A _5267_/A vssd1 vssd1 vccd1 vccd1
+ _5418_/B sky130_fd_sc_hd__mux4_1
XFILLER_114_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5348_ _7547_/Q _7437_/Q _7405_/Q _7389_/Q _5299_/A _4374_/A vssd1 vssd1 vccd1 vccd1
+ _5348_/X sky130_fd_sc_hd__mux4_1
Xoutput163 _5457_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[11] sky130_fd_sc_hd__buf_2
Xoutput185 _5491_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[31] sky130_fd_sc_hd__buf_2
Xoutput174 _5479_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5279_ _5279_/A vssd1 vssd1 vccd1 vccd1 _5279_/X sky130_fd_sc_hd__clkbuf_1
X_7018_ _6919_/A _6450_/A _7024_/S vssd1 vssd1 vccd1 vccd1 _7019_/B sky130_fd_sc_hd__mux2_1
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3077_ _6262_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3077_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6038__320 _6041__323/A vssd1 vssd1 vccd1 vccd1 _7246_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2627_ clkbuf_0__2627_/X vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4650_ _4249_/X _7238_/Q _4652_/S vssd1 vssd1 vccd1 vccd1 _4651_/A sky130_fd_sc_hd__mux2_1
Xinput21 caravel_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_2
Xinput10 caravel_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_4
X_3601_ _7700_/Q _3600_/X _3604_/S vssd1 vssd1 vccd1 vccd1 _3602_/A sky130_fd_sc_hd__mux2_1
Xinput32 caravel_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_4
X_6320_ _6320_/A vssd1 vssd1 vccd1 vccd1 _6320_/X sky130_fd_sc_hd__buf_1
X_4581_ _4581_/A vssd1 vssd1 vccd1 vccd1 _4581_/X sky130_fd_sc_hd__buf_2
Xinput54 wbs_data_i[0] vssd1 vssd1 vccd1 vccd1 _6908_/A sky130_fd_sc_hd__buf_12
Xinput43 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _5591_/B sky130_fd_sc_hd__clkbuf_2
X_3532_ _3532_/A vssd1 vssd1 vccd1 vccd1 _7711_/D sky130_fd_sc_hd__clkbuf_1
Xinput87 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _5748_/A sky130_fd_sc_hd__buf_6
Xinput65 wbs_data_i[1] vssd1 vssd1 vccd1 vccd1 _4976_/A sky130_fd_sc_hd__clkbuf_4
Xinput76 wbs_data_i[2] vssd1 vssd1 vccd1 vccd1 _3577_/A sky130_fd_sc_hd__buf_2
X_5202_ _7684_/Q _7607_/Q _5391_/S vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5133_ _7347_/Q vssd1 vssd1 vccd1 vccd1 _5270_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5064_ _5064_/A _5068_/B vssd1 vssd1 vccd1 vccd1 _5065_/A sky130_fd_sc_hd__and2_1
XFILLER_38_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4015_ _7490_/Q _3597_/X _4019_/S vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _5966_/A _5966_/B vssd1 vssd1 vccd1 vccd1 _5966_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5897_ _7212_/Q _7038_/Q _7260_/Q _7252_/Q _5818_/X _5819_/X vssd1 vssd1 vccd1 vccd1
+ _5897_/X sky130_fd_sc_hd__mux4_1
X_7705_ _7705_/CLK _7705_/D vssd1 vssd1 vccd1 vccd1 _7705_/Q sky130_fd_sc_hd__dfxtp_1
X_4917_ _4917_/A vssd1 vssd1 vccd1 vccd1 _7053_/D sky130_fd_sc_hd__clkbuf_1
X_7636_ _7636_/CLK _7636_/D vssd1 vssd1 vccd1 vccd1 _7636_/Q sky130_fd_sc_hd__dfxtp_1
X_4848_ _4820_/X _7121_/Q _4856_/S vssd1 vssd1 vccd1 vccd1 _4849_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2715_ _5694_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2715_/X sky130_fd_sc_hd__clkbuf_16
X_7567_ _7567_/CLK _7567_/D vssd1 vssd1 vccd1 vccd1 _7567_/Q sky130_fd_sc_hd__dfxtp_1
X_4779_ _4779_/A vssd1 vssd1 vccd1 vccd1 _7148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7498_ _7652_/CLK _7498_/D vssd1 vssd1 vccd1 vccd1 _7498_/Q sky130_fd_sc_hd__dfxtp_1
X_6518_ _6579_/C _6599_/A _6518_/C vssd1 vssd1 vccd1 vccd1 _6519_/A sky130_fd_sc_hd__and3b_1
X_6449_ _6448_/B _6448_/C _7507_/Q vssd1 vssd1 vccd1 vccd1 _6454_/B sky130_fd_sc_hd__a21oi_1
XFILLER_106_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6341__471 _6342__472/A vssd1 vssd1 vccd1 vccd1 _7413_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6665__110 _6666__111/A vssd1 vssd1 vccd1 vccd1 _7554_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6383__505 _6387__509/A vssd1 vssd1 vccd1 vccd1 _7447_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5820_ _7448_/Q _7440_/Q _7424_/Q _7416_/Q _5818_/X _5819_/X vssd1 vssd1 vccd1 vccd1
+ _5821_/B sky130_fd_sc_hd__mux4_1
XFILLER_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5751_ _5751_/A vssd1 vssd1 vccd1 vccd1 _7186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4702_ _4569_/X _7183_/Q _4706_/S vssd1 vssd1 vccd1 vccd1 _4703_/A sky130_fd_sc_hd__mux2_1
X_7421_ _7421_/CLK _7421_/D vssd1 vssd1 vccd1 vccd1 _7421_/Q sky130_fd_sc_hd__dfxtp_1
X_5682_ _5688_/A vssd1 vssd1 vccd1 vccd1 _5682_/X sky130_fd_sc_hd__buf_1
X_4633_ _4633_/A vssd1 vssd1 vccd1 vccd1 _7246_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4564_ _4560_/X _7273_/Q _4576_/S vssd1 vssd1 vccd1 vccd1 _4565_/A sky130_fd_sc_hd__mux2_1
X_7352_ _7352_/CLK _7352_/D vssd1 vssd1 vccd1 vccd1 _7352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7283_ _7283_/CLK _7283_/D vssd1 vssd1 vccd1 vccd1 _7283_/Q sky130_fd_sc_hd__dfxtp_1
X_3515_ _3822_/A _6233_/A vssd1 vssd1 vccd1 vccd1 _3711_/C sky130_fd_sc_hd__nor2_2
X_5661__223 _5661__223/A vssd1 vssd1 vccd1 vccd1 _7117_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4495_ _4495_/A vssd1 vssd1 vccd1 vccd1 _7307_/D sky130_fd_sc_hd__clkbuf_1
X_6234_ _7010_/A _6234_/B _6234_/C _6921_/C vssd1 vssd1 vccd1 vccd1 _6235_/A sky130_fd_sc_hd__and4_1
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6165_/A _6165_/B _6165_/C _6165_/D vssd1 vssd1 vccd1 vccd1 _6889_/A sky130_fd_sc_hd__or4_2
XFILLER_97_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _7731_/Q _7730_/Q _7729_/Q _7728_/Q vssd1 vssd1 vccd1 vccd1 _6450_/B sky130_fd_sc_hd__nor4_4
X_5116_ _7093_/Q _7094_/Q _7089_/Q _7090_/Q vssd1 vssd1 vccd1 vccd1 _5118_/B sky130_fd_sc_hd__or4_1
X_5047_ _5047_/A vssd1 vssd1 vccd1 vccd1 _5047_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6284__425 _6288__429/A vssd1 vssd1 vccd1 vccd1 _7367_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6998_ _6981_/X _6998_/B vssd1 vssd1 vccd1 vccd1 _6999_/A sky130_fd_sc_hd__and2b_1
X_5949_ _5888_/A _5948_/X _5929_/X vssd1 vssd1 vccd1 vccd1 _5949_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7619_ _7619_/CLK _7619_/D vssd1 vssd1 vccd1 vccd1 _7619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2629_ _5505_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2629_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2961_ clkbuf_0__2961_/X vssd1 vssd1 vccd1 vccd1 _6065__342/A sky130_fd_sc_hd__clkbuf_16
X_6729__162 _6729__162/A vssd1 vssd1 vccd1 vccd1 _7606_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4280_ _4280_/A vssd1 vssd1 vccd1 vccd1 _7385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6348__477 _6350__479/A vssd1 vssd1 vccd1 vccd1 _7419_/CLK sky130_fd_sc_hd__inv_2
X_6921_ _6921_/A _6921_/B _6921_/C vssd1 vssd1 vccd1 vccd1 _6922_/A sky130_fd_sc_hd__and3_1
X_6852_ _7650_/Q vssd1 vssd1 vccd1 vccd1 _6863_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3995_ _3995_/A vssd1 vssd1 vccd1 vccd1 _7520_/D sky130_fd_sc_hd__clkbuf_1
X_6783_ _6784_/A _6821_/A vssd1 vssd1 vccd1 vccd1 _6783_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4616_ _7253_/Q _3914_/A _4616_/S vssd1 vssd1 vccd1 vccd1 _4617_/A sky130_fd_sc_hd__mux2_1
X_7404_ _7404_/CLK _7404_/D vssd1 vssd1 vccd1 vccd1 _7404_/Q sky130_fd_sc_hd__dfxtp_1
X_5596_ _7082_/Q _5053_/A _5602_/S vssd1 vssd1 vccd1 vccd1 _5597_/A sky130_fd_sc_hd__mux2_1
X_7335_ _7335_/CLK _7335_/D vssd1 vssd1 vccd1 vccd1 _7335_/Q sky130_fd_sc_hd__dfxtp_1
X_4547_ _4547_/A vssd1 vssd1 vccd1 vccd1 _7283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7266_ _7266_/CLK _7266_/D vssd1 vssd1 vccd1 vccd1 _7266_/Q sky130_fd_sc_hd__dfxtp_1
X_4478_ _5888_/A _4482_/A vssd1 vssd1 vccd1 vccd1 _4479_/B sky130_fd_sc_hd__or2_1
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6251__402 _6252__403/A vssd1 vssd1 vccd1 vccd1 _7342_/CLK sky130_fd_sc_hd__inv_2
X_6217_ _6217_/A vssd1 vssd1 vccd1 vccd1 _7321_/D sky130_fd_sc_hd__clkbuf_1
X_7197_ _7727_/CLK _7197_/D vssd1 vssd1 vccd1 vccd1 _7197_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6148_ _6777_/A _6789_/A _6143_/Y _6788_/A _6147_/Y vssd1 vssd1 vccd1 vccd1 _6157_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_23 _7553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5522__193 _5522__193/A vssd1 vssd1 vccd1 vccd1 _7050_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_34 _5049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_12 _4340_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_45 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_56 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_67 _5492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_89 _7545_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_78 _5555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5668__229 _5668__229/A vssd1 vssd1 vccd1 vccd1 _7123_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3091_ clkbuf_0__3091_/X vssd1 vssd1 vccd1 vccd1 _6338__469/A sky130_fd_sc_hd__clkbuf_16
XFILLER_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6191__371 _6191__371/A vssd1 vssd1 vccd1 vccd1 _7301_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3780_ _3735_/X _7604_/Q _3786_/S vssd1 vssd1 vccd1 vccd1 _3781_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__3289_ clkbuf_0__3289_/X vssd1 vssd1 vccd1 vccd1 _6743__174/A sky130_fd_sc_hd__clkbuf_16
X_5450_ _5450_/A vssd1 vssd1 vccd1 vccd1 _5450_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4401_ _4416_/S vssd1 vssd1 vccd1 vccd1 _4410_/S sky130_fd_sc_hd__clkbuf_2
X_5381_ _5381_/A _5381_/B vssd1 vssd1 vccd1 vccd1 _5381_/Y sky130_fd_sc_hd__nor2_1
X_6710__147 _6710__147/A vssd1 vssd1 vccd1 vccd1 _7591_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7120_ _7120_/CLK _7120_/D vssd1 vssd1 vccd1 vccd1 _7120_/Q sky130_fd_sc_hd__dfxtp_1
X_4332_ _7364_/Q _4331_/X _4335_/S vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4263_ _4263_/A vssd1 vssd1 vccd1 vccd1 _7392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7051_ _7051_/CLK _7051_/D vssd1 vssd1 vccd1 vccd1 _7051_/Q sky130_fd_sc_hd__dfxtp_1
X_6002_ _7399_/Q _7241_/Q _7557_/Q _7463_/Q _5925_/A _5861_/X vssd1 vssd1 vccd1 vccd1
+ _6003_/B sky130_fd_sc_hd__mux4_1
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4194_ _4209_/S vssd1 vssd1 vccd1 vccd1 _4203_/S sky130_fd_sc_hd__buf_2
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6904_ _7665_/Q _6893_/B _6903_/X _6886_/X vssd1 vssd1 vccd1 vccd1 _7665_/D sky130_fd_sc_hd__o211a_1
XFILLER_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6966__52 _6968__54/A vssd1 vssd1 vccd1 vccd1 _7708_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6835_ _7646_/Q _6835_/B vssd1 vssd1 vccd1 vccd1 _6836_/B sky130_fd_sc_hd__or2_1
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6396__515 _6400__519/A vssd1 vssd1 vccd1 vccd1 _7457_/CLK sky130_fd_sc_hd__inv_2
X_3978_ _3978_/A vssd1 vssd1 vccd1 vccd1 _7528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5579_ _5706_/A vssd1 vssd1 vccd1 vccd1 _5579_/X sky130_fd_sc_hd__buf_1
X_7318_ _7318_/CLK _7318_/D vssd1 vssd1 vccd1 vccd1 _7318_/Q sky130_fd_sc_hd__dfxtp_1
X_7249_ _7249_/CLK _7249_/D vssd1 vssd1 vccd1 vccd1 _7249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6032__315 _6036__319/A vssd1 vssd1 vccd1 vccd1 _7241_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6297__435 _6298__436/A vssd1 vssd1 vccd1 vccd1 _7377_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__3074_ clkbuf_0__3074_/X vssd1 vssd1 vccd1 vccd1 _6256__406/A sky130_fd_sc_hd__clkbuf_16
X_6258__408 _6259__409/A vssd1 vssd1 vccd1 vccd1 _7348_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5529__199 _5529__199/A vssd1 vssd1 vccd1 vccd1 _7056_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput8 caravel_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4950_ _3816_/X _7037_/Q _4952_/S vssd1 vssd1 vccd1 vccd1 _4951_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3901_ _4121_/A _4642_/B vssd1 vssd1 vccd1 vccd1 _3924_/S sky130_fd_sc_hd__or2_2
XFILLER_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4881_ _4881_/A vssd1 vssd1 vccd1 vccd1 _7106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3832_ _3741_/X _7586_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3833_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6551_ _6553_/B _6556_/B _6562_/C vssd1 vssd1 vccd1 vccd1 _6551_/X sky130_fd_sc_hd__and3_1
X_3763_ _3763_/A vssd1 vssd1 vccd1 vccd1 _7612_/D sky130_fd_sc_hd__clkbuf_1
X_3694_ _3694_/A vssd1 vssd1 vccd1 vccd1 _7637_/D sky130_fd_sc_hd__clkbuf_1
X_6198__377 _6199__378/A vssd1 vssd1 vccd1 vccd1 _7307_/CLK sky130_fd_sc_hd__inv_2
X_6482_ _6483_/A _6483_/B _6483_/C _6483_/D vssd1 vssd1 vccd1 vccd1 _6482_/X sky130_fd_sc_hd__a31o_1
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5433_ _5433_/A _5433_/B _5433_/C vssd1 vssd1 vccd1 vccd1 _5433_/X sky130_fd_sc_hd__or3_1
X_5364_ _7522_/Q _7143_/Q _5403_/S vssd1 vssd1 vccd1 vccd1 _5364_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4315_ _4315_/A vssd1 vssd1 vccd1 vccd1 _7370_/D sky130_fd_sc_hd__clkbuf_1
X_7103_ _5496_/A _7103_/D vssd1 vssd1 vccd1 vccd1 _7103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5295_ _5349_/S _5294_/X _5178_/A vssd1 vssd1 vccd1 vccd1 _5295_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4246_ _7672_/Q vssd1 vssd1 vccd1 vccd1 _4246_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3093_ _6345_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3093_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7034_ _7034_/A _7034_/B vssd1 vssd1 vccd1 vccd1 _7035_/A sky130_fd_sc_hd__or2_1
X_4177_ _4094_/X _7423_/Q _4185_/S vssd1 vssd1 vccd1 vccd1 _4178_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6404__522 _6406__524/A vssd1 vssd1 vccd1 vccd1 _7464_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6818_ _6818_/A vssd1 vssd1 vccd1 vccd1 _7642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2712_ clkbuf_0__2712_/X vssd1 vssd1 vccd1 vccd1 _5681__239/A sky130_fd_sc_hd__clkbuf_16
XFILLER_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6305__442 _6307__444/A vssd1 vssd1 vccd1 vccd1 _7384_/CLK sky130_fd_sc_hd__inv_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3271_ clkbuf_0__3271_/X vssd1 vssd1 vccd1 vccd1 _6650__99/A sky130_fd_sc_hd__clkbuf_16
X_6960__47 _6961__48/A vssd1 vssd1 vccd1 vccd1 _7703_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__3057_ clkbuf_0__3057_/X vssd1 vssd1 vccd1 vccd1 _6214_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6078__348 _6079__349/A vssd1 vssd1 vccd1 vccd1 _7277_/CLK sky130_fd_sc_hd__inv_2
X_5080_ _5080_/A vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4100_ _7673_/Q vssd1 vssd1 vccd1 vccd1 _4100_/X sky130_fd_sc_hd__clkbuf_2
X_4031_ _3914_/X _7483_/Q _4031_/S vssd1 vssd1 vccd1 vccd1 _4032_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5982_ _7398_/Q _7240_/Q _7556_/Q _7462_/Q _5925_/A _4468_/A vssd1 vssd1 vccd1 vccd1
+ _5983_/B sky130_fd_sc_hd__mux4_1
XFILLER_92_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4933_ _4933_/A vssd1 vssd1 vccd1 vccd1 _7046_/D sky130_fd_sc_hd__clkbuf_1
X_7721_ _7722_/CLK _7721_/D vssd1 vssd1 vccd1 vccd1 _7721_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7652_ _7652_/CLK _7652_/D vssd1 vssd1 vccd1 vccd1 _7652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4864_ _4864_/A _4864_/B vssd1 vssd1 vccd1 vccd1 _4880_/S sky130_fd_sc_hd__or2_2
X_3815_ _3815_/A vssd1 vssd1 vccd1 vccd1 _7592_/D sky130_fd_sc_hd__clkbuf_1
X_7583_ _7583_/CLK _7583_/D vssd1 vssd1 vccd1 vccd1 _7583_/Q sky130_fd_sc_hd__dfxtp_1
X_6206__384 _6206__384/A vssd1 vssd1 vccd1 vccd1 _7314_/CLK sky130_fd_sc_hd__inv_2
X_4795_ _4795_/A vssd1 vssd1 vccd1 vccd1 _7141_/D sky130_fd_sc_hd__clkbuf_1
X_6603_ _6601_/Y _6599_/C _6602_/X _6569_/A vssd1 vssd1 vccd1 vccd1 _7512_/D sky130_fd_sc_hd__o211a_1
X_3746_ _3746_/A vssd1 vssd1 vccd1 vccd1 _7617_/D sky130_fd_sc_hd__clkbuf_1
X_6534_ _6534_/A vssd1 vssd1 vccd1 vccd1 _6583_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6465_ _6158_/A _6112_/A _6464_/Y vssd1 vssd1 vccd1 vccd1 _6500_/B sky130_fd_sc_hd__a21o_1
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3677_ _3677_/A vssd1 vssd1 vccd1 vccd1 _7681_/D sky130_fd_sc_hd__clkbuf_1
X_5416_ _7293_/Q _7079_/Q _7706_/Q _7367_/Q _5303_/X _5299_/X vssd1 vssd1 vccd1 vccd1
+ _5416_/X sky130_fd_sc_hd__mux4_1
Xoutput142 _5039_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[28] sky130_fd_sc_hd__buf_2
Xoutput120 _5067_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[9] sky130_fd_sc_hd__buf_2
Xoutput131 _5017_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[18] sky130_fd_sc_hd__buf_2
Xoutput153 _4996_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[9] sky130_fd_sc_hd__buf_2
X_5347_ _7135_/Q _7058_/Q _7050_/Q _7271_/Q _5267_/A _4381_/A vssd1 vssd1 vccd1 vccd1
+ _5347_/X sky130_fd_sc_hd__mux4_1
Xoutput164 _5460_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[12] sky130_fd_sc_hd__buf_2
Xoutput175 _5480_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput186 _5312_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_99_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5278_ _5278_/A _5278_/B vssd1 vssd1 vccd1 vccd1 _5279_/A sky130_fd_sc_hd__or2_1
X_4229_ _4578_/A vssd1 vssd1 vccd1 vccd1 _4229_/X sky130_fd_sc_hd__buf_2
X_7017_ _7017_/A vssd1 vssd1 vccd1 vccd1 _7726_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3076_ _6261_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3076_/X sky130_fd_sc_hd__clkbuf_16
X_6723__157 _6724__158/A vssd1 vssd1 vccd1 vccd1 _7601_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2626_ clkbuf_0__2626_/X vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6933__25 _6934__26/A vssd1 vssd1 vccd1 vccd1 _7681_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 caravel_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_2
Xinput11 caravel_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_4
X_4580_ _4580_/A vssd1 vssd1 vccd1 vccd1 _7268_/D sky130_fd_sc_hd__clkbuf_1
X_3600_ _7322_/Q vssd1 vssd1 vccd1 vccd1 _3600_/X sky130_fd_sc_hd__buf_4
Xinput33 caravel_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__3109_ clkbuf_0__3109_/X vssd1 vssd1 vccd1 vccd1 _6424__57/A sky130_fd_sc_hd__clkbuf_16
X_3531_ _3530_/X _7711_/Q _3535_/S vssd1 vssd1 vccd1 vccd1 _3532_/A sky130_fd_sc_hd__mux2_1
Xinput44 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _5049_/A sky130_fd_sc_hd__buf_4
Xinput55 wbs_data_i[10] vssd1 vssd1 vccd1 vccd1 _4997_/A sky130_fd_sc_hd__buf_4
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput88 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _5766_/A sky130_fd_sc_hd__buf_8
Xinput66 wbs_data_i[20] vssd1 vssd1 vccd1 vccd1 _5020_/A sky130_fd_sc_hd__buf_4
Xinput77 wbs_data_i[30] vssd1 vssd1 vccd1 vccd1 _5042_/A sky130_fd_sc_hd__buf_4
XFILLER_6_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5201_ _4375_/A _5201_/B vssd1 vssd1 vccd1 vccd1 _5201_/X sky130_fd_sc_hd__and2b_1
X_5132_ _5303_/A vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__buf_2
XFILLER_111_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5063_ _5063_/A vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__clkbuf_1
X_4014_ _4014_/A vssd1 vssd1 vccd1 vccd1 _7491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5965_ _7627_/Q _7619_/Q _7603_/Q _7595_/Q _5823_/X _5925_/X vssd1 vssd1 vccd1 vccd1
+ _5966_/B sky130_fd_sc_hd__mux4_2
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5896_ _5894_/X _5895_/X _5959_/S vssd1 vssd1 vccd1 vccd1 _5896_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7704_ _7704_/CLK _7704_/D vssd1 vssd1 vccd1 vccd1 _7704_/Q sky130_fd_sc_hd__dfxtp_1
X_4916_ _4843_/X _7053_/Q _4916_/S vssd1 vssd1 vccd1 vccd1 _4917_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7635_ _7635_/CLK _7635_/D vssd1 vssd1 vccd1 vccd1 _7635_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2714_ _5688_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2714_/X sky130_fd_sc_hd__clkbuf_16
X_4847_ _4862_/S vssd1 vssd1 vccd1 vccd1 _4856_/S sky130_fd_sc_hd__buf_2
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7566_ _7566_/CLK _7566_/D vssd1 vssd1 vccd1 vccd1 _7566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4778_ _7148_/Q _4337_/X _4782_/S vssd1 vssd1 vccd1 vccd1 _4779_/A sky130_fd_sc_hd__mux2_1
X_3729_ _3729_/A vssd1 vssd1 vccd1 vccd1 _7622_/D sky130_fd_sc_hd__clkbuf_1
X_7497_ _7525_/CLK _7497_/D vssd1 vssd1 vccd1 vccd1 _7497_/Q sky130_fd_sc_hd__dfxtp_1
X_6517_ _6534_/A _6516_/X _6610_/B vssd1 vssd1 vccd1 vccd1 _6518_/C sky130_fd_sc_hd__o21ai_1
X_6448_ _7507_/Q _6448_/B _6448_/C vssd1 vssd1 vccd1 vccd1 _6454_/A sky130_fd_sc_hd__and3_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3059_ _6214_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3059_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5750_ _4993_/A _7186_/Q _5758_/S vssd1 vssd1 vccd1 vccd1 _5751_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4701_/A vssd1 vssd1 vccd1 vccd1 _7184_/D sky130_fd_sc_hd__clkbuf_1
X_4632_ _4249_/X _7246_/Q _4634_/S vssd1 vssd1 vccd1 vccd1 _4633_/A sky130_fd_sc_hd__mux2_1
X_7420_ _7420_/CLK _7420_/D vssd1 vssd1 vccd1 vccd1 _7420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4563_ _4585_/S vssd1 vssd1 vccd1 vccd1 _4576_/S sky130_fd_sc_hd__buf_2
X_7351_ _7351_/CLK _7351_/D vssd1 vssd1 vccd1 vccd1 _7351_/Q sky130_fd_sc_hd__dfxtp_2
X_7282_ _7282_/CLK _7282_/D vssd1 vssd1 vccd1 vccd1 _7282_/Q sky130_fd_sc_hd__dfxtp_1
X_6302_ _6308_/A vssd1 vssd1 vccd1 vccd1 _6302_/X sky130_fd_sc_hd__buf_1
X_4494_ _4220_/X _7307_/Q _4498_/S vssd1 vssd1 vccd1 vccd1 _4495_/A sky130_fd_sc_hd__mux2_1
X_3514_ _3610_/A _3513_/X _3611_/A vssd1 vssd1 vccd1 vccd1 _6233_/A sky130_fd_sc_hd__a21o_4
X_6233_ _6233_/A _6233_/B vssd1 vssd1 vccd1 vccd1 _6921_/C sky130_fd_sc_hd__nor2_4
Xclkbuf_1_0__f__3099_ clkbuf_0__3099_/X vssd1 vssd1 vccd1 vccd1 _6379__502/A sky130_fd_sc_hd__clkbuf_16
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6771_/B _6774_/B _6164_/C vssd1 vssd1 vccd1 vccd1 _6165_/D sky130_fd_sc_hd__or3_1
XFILLER_111_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6492_/B vssd1 vssd1 vccd1 vccd1 _6163_/A sky130_fd_sc_hd__clkbuf_2
X_5115_ _7095_/Q _7096_/Q _5645_/B _5115_/D vssd1 vssd1 vccd1 vccd1 _5118_/A sky130_fd_sc_hd__or4_1
X_5046_ _5046_/A _5046_/B vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__and2_1
XFILLER_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6997_ _4999_/A _7721_/Q _7000_/S vssd1 vssd1 vccd1 vccd1 _6998_/B sky130_fd_sc_hd__mux2_1
XFILLER_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5948_ _7412_/Q _7380_/Q _7711_/Q _7634_/Q _5819_/X _5884_/X vssd1 vssd1 vccd1 vccd1
+ _5948_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5879_ _5865_/X _5878_/X _5833_/X vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__a21bo_1
X_7618_ _7618_/CLK _7618_/D vssd1 vssd1 vccd1 vccd1 _7618_/Q sky130_fd_sc_hd__dfxtp_1
X_7549_ _7549_/CLK _7549_/D vssd1 vssd1 vccd1 vccd1 _7549_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__2628_ _5499_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2628_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2960_ clkbuf_0__2960_/X vssd1 vssd1 vccd1 vccd1 _6061__339/A sky130_fd_sc_hd__clkbuf_16
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7723_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_71_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6920_ _6920_/A vssd1 vssd1 vccd1 vccd1 _7672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6851_ _6851_/A vssd1 vssd1 vccd1 vccd1 _7649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3994_ _3656_/X _7520_/Q _3994_/S vssd1 vssd1 vccd1 vccd1 _3995_/A sky130_fd_sc_hd__mux2_1
X_6782_ _7639_/Q vssd1 vssd1 vccd1 vccd1 _6794_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6760__12 _6761__13/A vssd1 vssd1 vccd1 vccd1 _7631_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4615_ _4615_/A vssd1 vssd1 vccd1 vccd1 _7254_/D sky130_fd_sc_hd__clkbuf_1
X_7403_ _7403_/CLK _7403_/D vssd1 vssd1 vccd1 vccd1 _7403_/Q sky130_fd_sc_hd__dfxtp_1
X_5595_ _5595_/A vssd1 vssd1 vccd1 vccd1 _7081_/D sky130_fd_sc_hd__clkbuf_1
X_4546_ _7283_/Q _3905_/A _4552_/S vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__mux2_1
X_7334_ _7334_/CLK _7334_/D vssd1 vssd1 vccd1 vccd1 _7334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7265_ _7265_/CLK _7265_/D vssd1 vssd1 vccd1 vccd1 _7265_/Q sky130_fd_sc_hd__dfxtp_1
X_4477_ _4477_/A _4477_/B vssd1 vssd1 vccd1 vccd1 _4482_/A sky130_fd_sc_hd__and2_1
X_6290__430 _6294__434/A vssd1 vssd1 vccd1 vccd1 _7372_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6216_ _7659_/Q _6220_/B vssd1 vssd1 vccd1 vccd1 _6217_/A sky130_fd_sc_hd__and2_1
X_7196_ _7670_/CLK _7196_/D vssd1 vssd1 vccd1 vccd1 _7196_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6147_ _6450_/B _6792_/C vssd1 vssd1 vccd1 vccd1 _6147_/Y sky130_fd_sc_hd__xnor2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_24 _7554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_13 _4343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_46 _4993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_68 _5895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_57 _3813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_35 _5049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5029_ _5029_/A _5035_/B vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__and2_1
XFILLER_72_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_79 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3090_ clkbuf_0__3090_/X vssd1 vssd1 vccd1 vccd1 _6331__463/A sky130_fd_sc_hd__clkbuf_16
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__3288_ clkbuf_0__3288_/X vssd1 vssd1 vccd1 vccd1 _6736__168/A sky130_fd_sc_hd__clkbuf_16
XFILLER_12_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ _4400_/A _4506_/B vssd1 vssd1 vccd1 vccd1 _4416_/S sky130_fd_sc_hd__nor2_2
X_6200__379 _6200__379/A vssd1 vssd1 vccd1 vccd1 _7309_/CLK sky130_fd_sc_hd__inv_2
X_5380_ _5380_/A _5380_/B _5380_/C _5587_/C vssd1 vssd1 vccd1 vccd1 _5381_/B sky130_fd_sc_hd__or4_1
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4331_ _7325_/Q vssd1 vssd1 vccd1 vccd1 _4331_/X sky130_fd_sc_hd__clkbuf_4
X_4262_ _4261_/X _7392_/Q _4262_/S vssd1 vssd1 vccd1 vccd1 _4263_/A sky130_fd_sc_hd__mux2_1
X_7050_ _7050_/CLK _7050_/D vssd1 vssd1 vccd1 vccd1 _7050_/Q sky130_fd_sc_hd__dfxtp_1
X_6354__482 _6355__483/A vssd1 vssd1 vccd1 vccd1 _7424_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6001_ _6001_/A _6001_/B vssd1 vssd1 vccd1 vccd1 _6001_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4193_ _4283_/A _4239_/A vssd1 vssd1 vccd1 vccd1 _4209_/S sky130_fd_sc_hd__or2_2
XFILLER_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6903_ _7666_/Q _6903_/B vssd1 vssd1 vccd1 vccd1 _6903_/X sky130_fd_sc_hd__or2_1
X_6678__121 _6681__124/A vssd1 vssd1 vccd1 vccd1 _7565_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__2962_ _6068_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2962_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6834_ _6847_/D vssd1 vssd1 vccd1 vccd1 _6843_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3977_ _3660_/X _7528_/Q _3981_/S vssd1 vssd1 vccd1 vccd1 _3978_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5647_ _5647_/A _5647_/B _5588_/X vssd1 vssd1 vccd1 vccd1 _7104_/D sky130_fd_sc_hd__nor3b_1
X_5708__260 _5712__264/A vssd1 vssd1 vccd1 vccd1 _7154_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7317_ _7317_/CLK _7317_/D vssd1 vssd1 vccd1 vccd1 _7317_/Q sky130_fd_sc_hd__dfxtp_1
X_4529_ _4529_/A vssd1 vssd1 vccd1 vccd1 _7292_/D sky130_fd_sc_hd__clkbuf_1
X_7248_ _7248_/CLK _7248_/D vssd1 vssd1 vccd1 vccd1 _7248_/Q sky130_fd_sc_hd__dfxtp_1
X_7179_ _7179_/CLK _7179_/D vssd1 vssd1 vccd1 vccd1 _7179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5674__234 _5674__234/A vssd1 vssd1 vccd1 vccd1 _7128_/CLK sky130_fd_sc_hd__inv_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__3073_ clkbuf_0__3073_/X vssd1 vssd1 vccd1 vccd1 _6253__404/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5802__292 _5804__294/A vssd1 vssd1 vccd1 vccd1 _7210_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 caravel_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3900_ _4095_/A _4095_/B _3900_/C vssd1 vssd1 vccd1 vccd1 _4642_/B sky130_fd_sc_hd__or3_4
X_4880_ _4843_/X _7106_/Q _4880_/S vssd1 vssd1 vccd1 vccd1 _4881_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3831_ _3831_/A vssd1 vssd1 vccd1 vccd1 _7587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3762_ _3644_/X _7612_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3763_/A sky130_fd_sc_hd__mux2_1
X_6550_ _6566_/A _6550_/B _6550_/C vssd1 vssd1 vccd1 vccd1 _6550_/X sky130_fd_sc_hd__and3_1
XFILLER_118_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3693_ _3469_/X _7637_/Q _3701_/S vssd1 vssd1 vccd1 vccd1 _3694_/A sky130_fd_sc_hd__mux2_1
X_6481_ _6481_/A _7505_/Q vssd1 vssd1 vccd1 vccd1 _6483_/D sky130_fd_sc_hd__xor2_1
XFILLER_118_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5432_ _5428_/X _5430_/X _5431_/X _5415_/A _4368_/A vssd1 vssd1 vccd1 vccd1 _5433_/C
+ sky130_fd_sc_hd__o221a_1
X_5363_ _5363_/A _5363_/B vssd1 vssd1 vccd1 vccd1 _5363_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4314_ _4229_/X _7370_/Q _4318_/S vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__mux2_1
X_7102_ _7727_/CLK _7102_/D vssd1 vssd1 vccd1 vccd1 _7102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5294_ _7173_/Q _7305_/Q _7491_/Q _7181_/Q _5267_/A _5290_/S vssd1 vssd1 vccd1 vccd1
+ _5294_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_0__3092_ _6339_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3092_/X sky130_fd_sc_hd__clkbuf_16
X_4245_ _4245_/A vssd1 vssd1 vccd1 vccd1 _7398_/D sky130_fd_sc_hd__clkbuf_1
X_7033_ _6908_/A _7732_/Q _7033_/S vssd1 vssd1 vccd1 vccd1 _7034_/B sky130_fd_sc_hd__mux2_1
X_4176_ _4191_/S vssd1 vssd1 vccd1 vccd1 _4185_/S sky130_fd_sc_hd__buf_2
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6817_ _6821_/B _6817_/B _6872_/B vssd1 vssd1 vccd1 vccd1 _6818_/A sky130_fd_sc_hd__and3b_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2711_ clkbuf_0__2711_/X vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_74_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__3270_ clkbuf_0__3270_/X vssd1 vssd1 vccd1 vccd1 _6642__92/A sky130_fd_sc_hd__clkbuf_16
XFILLER_115_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3056_ clkbuf_0__3056_/X vssd1 vssd1 vccd1 vccd1 _6206__384/A sky130_fd_sc_hd__clkbuf_16
XFILLER_10_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6271__417 _6276__419/A vssd1 vssd1 vccd1 vccd1 _7357_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4030_ _4030_/A vssd1 vssd1 vccd1 vccd1 _7484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6618__74 _6618__74/A vssd1 vssd1 vccd1 vccd1 _7517_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5981_ _6001_/A _5981_/B vssd1 vssd1 vccd1 vccd1 _5981_/Y sky130_fd_sc_hd__nor2_1
X_4932_ _7046_/Q _4581_/A _4934_/S vssd1 vssd1 vccd1 vccd1 _4933_/A sky130_fd_sc_hd__mux2_1
X_7720_ _7722_/CLK _7720_/D vssd1 vssd1 vccd1 vccd1 _7720_/Q sky130_fd_sc_hd__dfxtp_4
X_7651_ _7655_/CLK _7651_/D vssd1 vssd1 vccd1 vccd1 _7651_/Q sky130_fd_sc_hd__dfxtp_1
X_4863_ _4863_/A vssd1 vssd1 vccd1 vccd1 _7114_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6602_ _7511_/Q _6566_/A _6604_/C _7512_/Q vssd1 vssd1 vccd1 vccd1 _6602_/X sky130_fd_sc_hd__a31o_1
XFILLER_119_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3814_ _7592_/Q _3813_/X _3820_/S vssd1 vssd1 vccd1 vccd1 _3815_/A sky130_fd_sc_hd__mux2_1
X_7582_ _7582_/CLK _7582_/D vssd1 vssd1 vccd1 vccd1 _7582_/Q sky130_fd_sc_hd__dfxtp_1
X_4794_ _7141_/Q _4575_/A _4794_/S vssd1 vssd1 vccd1 vccd1 _4795_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3745_ _3744_/X _7617_/Q _3745_/S vssd1 vssd1 vccd1 vccd1 _3746_/A sky130_fd_sc_hd__mux2_1
X_6533_ _6541_/C _6532_/C _6541_/B vssd1 vssd1 vccd1 vccd1 _6535_/B sky130_fd_sc_hd__a21o_1
XFILLER_118_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5809__298 _5810__299/A vssd1 vssd1 vccd1 vccd1 _7216_/CLK sky130_fd_sc_hd__inv_2
X_6464_ _7513_/Q vssd1 vssd1 vccd1 vccd1 _6464_/Y sky130_fd_sc_hd__inv_2
Xoutput110 _5103_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[25] sky130_fd_sc_hd__buf_2
XFILLER_118_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3676_ _3522_/X _7681_/Q _3682_/S vssd1 vssd1 vccd1 vccd1 _3677_/A sky130_fd_sc_hd__mux2_1
X_5415_ _5415_/A _5415_/B vssd1 vssd1 vccd1 vccd1 _5415_/X sky130_fd_sc_hd__or2_1
Xoutput143 _5041_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[29] sky130_fd_sc_hd__buf_2
Xoutput132 _5019_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput121 _4966_/B vssd1 vssd1 vccd1 vccd1 caravel_wb_cyc_o sky130_fd_sc_hd__buf_2
X_6395_ _6395_/A vssd1 vssd1 vccd1 vccd1 _6395_/X sky130_fd_sc_hd__buf_1
Xoutput154 _4965_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[0] sky130_fd_sc_hd__buf_2
XFILLER_99_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput165 _5463_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput176 _5483_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5346_ _6149_/A vssd1 vssd1 vccd1 vccd1 _6450_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput187 _5343_/Y vssd1 vssd1 vccd1 vccd1 wbs_data_o[4] sky130_fd_sc_hd__buf_2
X_5277_ _6119_/B _5236_/X _5275_/Y _5276_/X _5112_/X vssd1 vssd1 vccd1 vccd1 _5278_/B
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__3075_ _6260_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3075_/X sky130_fd_sc_hd__clkbuf_16
X_4228_ _4228_/A vssd1 vssd1 vccd1 vccd1 _7403_/D sky130_fd_sc_hd__clkbuf_1
X_7016_ _7031_/A _7016_/B vssd1 vssd1 vccd1 vccd1 _7017_/A sky130_fd_sc_hd__or2_1
X_6213__389 _6213__389/A vssd1 vssd1 vccd1 vccd1 _7319_/CLK sky130_fd_sc_hd__inv_2
X_4159_ _4094_/X _7431_/Q _4167_/S vssd1 vssd1 vccd1 vccd1 _4160_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6367__492 _6368__493/A vssd1 vssd1 vccd1 vccd1 _7434_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2625_ clkbuf_0__2625_/X vssd1 vssd1 vccd1 vccd1 _6260_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6084__353 _6085__354/A vssd1 vssd1 vccd1 vccd1 _7282_/CLK sky130_fd_sc_hd__inv_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6045__326 _6048__329/A vssd1 vssd1 vccd1 vccd1 _7252_/CLK sky130_fd_sc_hd__inv_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5687__244 _5687__244/A vssd1 vssd1 vccd1 vccd1 _7138_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 caravel_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_2
Xinput23 caravel_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_2
Xinput34 caravel_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__3108_ clkbuf_0__3108_/X vssd1 vssd1 vccd1 vccd1 _6427_/A sky130_fd_sc_hd__clkbuf_16
X_3530_ _3911_/A vssd1 vssd1 vccd1 vccd1 _3530_/X sky130_fd_sc_hd__buf_2
Xinput45 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _5051_/A sky130_fd_sc_hd__buf_4
Xinput78 wbs_data_i[31] vssd1 vssd1 vccd1 vccd1 _5044_/A sky130_fd_sc_hd__buf_4
Xinput89 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _5784_/A sky130_fd_sc_hd__buf_6
Xinput56 wbs_data_i[11] vssd1 vssd1 vccd1 vccd1 _4999_/A sky130_fd_sc_hd__buf_4
Xinput67 wbs_data_i[21] vssd1 vssd1 vccd1 vccd1 _5022_/A sky130_fd_sc_hd__buf_4
X_5200_ _7115_/Q _7163_/Q _5391_/S vssd1 vssd1 vccd1 vccd1 _5201_/B sky130_fd_sc_hd__mux2_1
X_5131_ _5205_/A vssd1 vssd1 vccd1 vccd1 _5131_/X sky130_fd_sc_hd__clkbuf_2
X_5062_ _5062_/A _5068_/B vssd1 vssd1 vccd1 vccd1 _5063_/A sky130_fd_sc_hd__and2_1
XFILLER_57_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4013_ _7491_/Q _3594_/X _4013_/S vssd1 vssd1 vccd1 vccd1 _4014_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6767__18 _6925__19/A vssd1 vssd1 vccd1 vccd1 _7637_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5964_ _6003_/A _5964_/B vssd1 vssd1 vccd1 vccd1 _5964_/Y sky130_fd_sc_hd__nor2_1
X_7703_ _7703_/CLK _7703_/D vssd1 vssd1 vccd1 vccd1 _7703_/Q sky130_fd_sc_hd__dfxtp_1
X_5895_ _7584_/Q _7576_/Q _7568_/Q _7482_/Q _5818_/X _4462_/A vssd1 vssd1 vccd1 vccd1
+ _5895_/X sky130_fd_sc_hd__mux4_2
XFILLER_80_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4915_ _4915_/A vssd1 vssd1 vccd1 vccd1 _7054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7634_ _7634_/CLK _7634_/D vssd1 vssd1 vccd1 vccd1 _7634_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2713_ _5682_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2713_/X sky130_fd_sc_hd__clkbuf_16
X_4846_ _4846_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4862_/S sky130_fd_sc_hd__or2_2
X_7565_ _7565_/CLK _7565_/D vssd1 vssd1 vccd1 vccd1 _7565_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ _4777_/A vssd1 vssd1 vccd1 vccd1 _7149_/D sky130_fd_sc_hd__clkbuf_1
X_6516_ _6236_/C _6510_/X _6515_/X _7497_/Q vssd1 vssd1 vccd1 vccd1 _6516_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3728_ _3546_/X _7622_/Q _3728_/S vssd1 vssd1 vccd1 vccd1 _3729_/A sky130_fd_sc_hd__mux2_1
X_7496_ _7510_/CLK _7496_/D vssd1 vssd1 vccd1 vccd1 _7496_/Q sky130_fd_sc_hd__dfxtp_1
X_3659_ _7323_/Q vssd1 vssd1 vccd1 vccd1 _4578_/A sky130_fd_sc_hd__buf_2
X_6447_ _6137_/A _6159_/A _6446_/B _6129_/A vssd1 vssd1 vccd1 vccd1 _6448_/C sky130_fd_sc_hd__o31ai_1
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5329_ _5315_/A _5324_/Y _5326_/X _5328_/Y vssd1 vssd1 vccd1 vccd1 _5337_/B sky130_fd_sc_hd__a31o_1
XFILLER_102_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3058_ _6208_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3058_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_90_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6417__533 _6418__534/A vssd1 vssd1 vccd1 vccd1 _7475_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4566_/X _7184_/Q _4706_/S vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4631_ _4631_/A vssd1 vssd1 vccd1 vccd1 _7247_/D sky130_fd_sc_hd__clkbuf_1
X_6672__116 _6675__119/A vssd1 vssd1 vccd1 vccd1 _7560_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4562_ _4562_/A _4918_/B vssd1 vssd1 vccd1 vccd1 _4585_/S sky130_fd_sc_hd__or2_1
XFILLER_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7350_ _7350_/CLK _7350_/D vssd1 vssd1 vccd1 vccd1 _7350_/Q sky130_fd_sc_hd__dfxtp_2
X_7281_ _7281_/CLK _7281_/D vssd1 vssd1 vccd1 vccd1 _7281_/Q sky130_fd_sc_hd__dfxtp_1
X_4493_ _4493_/A vssd1 vssd1 vccd1 vccd1 _7308_/D sky130_fd_sc_hd__clkbuf_1
X_3513_ _3513_/A vssd1 vssd1 vccd1 vccd1 _3513_/X sky130_fd_sc_hd__buf_4
X_6318__453 _6319__454/A vssd1 vssd1 vccd1 vccd1 _7395_/CLK sky130_fd_sc_hd__inv_2
X_6232_ _6232_/A vssd1 vssd1 vccd1 vccd1 _7328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5509__187 _5509__187/A vssd1 vssd1 vccd1 vccd1 _7043_/CLK sky130_fd_sc_hd__inv_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3098_ clkbuf_0__3098_/X vssd1 vssd1 vccd1 vccd1 _6373__497/A sky130_fd_sc_hd__clkbuf_16
X_6163_ _6163_/A _6791_/C vssd1 vssd1 vccd1 vccd1 _6164_/C sky130_fd_sc_hd__xnor2_1
XFILLER_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _7721_/Q _6446_/A _6127_/C _6093_/Y vssd1 vssd1 vccd1 vccd1 _6492_/B sky130_fd_sc_hd__or4b_2
X_5114_ _7097_/Q _7098_/Q _7099_/Q _7100_/Q vssd1 vssd1 vccd1 vccd1 _5115_/D sky130_fd_sc_hd__or4_1
X_5045_ _5045_/A vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6996_ _6996_/A vssd1 vssd1 vccd1 vccd1 _7720_/D sky130_fd_sc_hd__clkbuf_1
X_5947_ _5966_/A _5947_/B vssd1 vssd1 vccd1 vccd1 _5947_/Y sky130_fd_sc_hd__nor2_1
X_7617_ _7617_/CLK _7617_/D vssd1 vssd1 vccd1 vccd1 _7617_/Q sky130_fd_sc_hd__dfxtp_1
X_5878_ _3485_/Y _5868_/X _5872_/X _5876_/X _5882_/A vssd1 vssd1 vccd1 vccd1 _5878_/X
+ sky130_fd_sc_hd__a311o_1
X_4829_ _4828_/X _7127_/Q _4835_/S vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2627_ _5498_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2627_/X sky130_fd_sc_hd__clkbuf_16
X_7548_ _7548_/CLK _7548_/D vssd1 vssd1 vccd1 vccd1 _7548_/Q sky130_fd_sc_hd__dfxtp_1
X_7479_ _7479_/CLK _7479_/D vssd1 vssd1 vccd1 vccd1 _7479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5534__203 _5572__204/A vssd1 vssd1 vccd1 vccd1 _7060_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6736__168 _6736__168/A vssd1 vssd1 vccd1 vccd1 _7612_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6850_ _6857_/C _6850_/B _6859_/C vssd1 vssd1 vccd1 vccd1 _6851_/A sky130_fd_sc_hd__and3b_1
XFILLER_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6781_ _6781_/A vssd1 vssd1 vccd1 vccd1 _6781_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5801_ _5801_/A vssd1 vssd1 vccd1 vccd1 _7209_/D sky130_fd_sc_hd__clkbuf_1
X_3993_ _3993_/A vssd1 vssd1 vccd1 vccd1 _7521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5663_ _5663_/A vssd1 vssd1 vccd1 vccd1 _5663_/X sky130_fd_sc_hd__buf_1
X_4614_ _7254_/Q _3911_/A _4616_/S vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__mux2_1
X_7402_ _7402_/CLK _7402_/D vssd1 vssd1 vccd1 vccd1 _7402_/Q sky130_fd_sc_hd__dfxtp_2
X_5594_ _7081_/Q _5051_/A _5602_/S vssd1 vssd1 vccd1 vccd1 _5595_/A sky130_fd_sc_hd__mux2_1
X_4545_ _4545_/A vssd1 vssd1 vccd1 vccd1 _7284_/D sky130_fd_sc_hd__clkbuf_1
X_7333_ _7333_/CLK _7333_/D vssd1 vssd1 vccd1 vccd1 _7333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6058__336 _6061__339/A vssd1 vssd1 vccd1 vccd1 _7262_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7264_ _7264_/CLK _7264_/D vssd1 vssd1 vccd1 vccd1 _7264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4476_ _5899_/S vssd1 vssd1 vccd1 vccd1 _5888_/A sky130_fd_sc_hd__clkbuf_2
X_7195_ _7670_/CLK _7195_/D vssd1 vssd1 vccd1 vccd1 _7195_/Q sky130_fd_sc_hd__dfxtp_4
X_6146_ _6149_/A _7644_/Q vssd1 vssd1 vccd1 vccd1 _6792_/C sky130_fd_sc_hd__xnor2_2
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_14 _5106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_25 _7556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_47 _4995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_58 _3813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_36 _5049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6077_ _6077_/A vssd1 vssd1 vccd1 vccd1 _7276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5028_ _5028_/A vssd1 vssd1 vccd1 vccd1 _5028_/X sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_69 _5937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6979_ _5590_/A _6979_/B vssd1 vssd1 vccd1 vccd1 _6980_/A sky130_fd_sc_hd__and2b_1
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3287_ clkbuf_0__3287_/X vssd1 vssd1 vccd1 vccd1 _6729__162/A sky130_fd_sc_hd__clkbuf_16
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4330_ _4330_/A vssd1 vssd1 vccd1 vccd1 _7365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4261_ _7667_/Q vssd1 vssd1 vccd1 vccd1 _4261_/X sky130_fd_sc_hd__buf_2
XFILLER_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6000_ _7455_/Q _7447_/Q _7431_/Q _7423_/Q _5851_/X _5852_/X vssd1 vssd1 vccd1 vccd1
+ _6001_/B sky130_fd_sc_hd__mux4_1
X_4192_ _4192_/A vssd1 vssd1 vccd1 vccd1 _7416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2961_ _6062_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2961_/X sky130_fd_sc_hd__clkbuf_16
X_6902_ _7665_/Q _6892_/X _6901_/X _6886_/X vssd1 vssd1 vccd1 vccd1 _7664_/D sky130_fd_sc_hd__o211a_1
X_6833_ _7646_/Q _7645_/Q _6833_/C _6833_/D vssd1 vssd1 vccd1 vccd1 _6847_/D sky130_fd_sc_hd__and4_1
Xclkbuf_1_0__f__2719_ clkbuf_0__2719_/X vssd1 vssd1 vccd1 vccd1 _5718__269/A sky130_fd_sc_hd__clkbuf_16
XFILLER_35_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6361__487 _6363__489/A vssd1 vssd1 vccd1 vccd1 _7429_/CLK sky130_fd_sc_hd__inv_2
X_3976_ _3976_/A vssd1 vssd1 vccd1 vccd1 _7529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6695_ _6701_/A vssd1 vssd1 vccd1 vccd1 _6695_/X sky130_fd_sc_hd__buf_1
X_5646_ _5587_/B _5380_/C _5645_/Y _7034_/A vssd1 vssd1 vccd1 vccd1 _5647_/A sky130_fd_sc_hd__a31o_1
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7316_ _7316_/CLK _7316_/D vssd1 vssd1 vccd1 vccd1 _7316_/Q sky130_fd_sc_hd__dfxtp_2
X_4528_ _4217_/X _7292_/Q _4534_/S vssd1 vssd1 vccd1 vccd1 _4529_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7247_ _7247_/CLK _7247_/D vssd1 vssd1 vccd1 vccd1 _7247_/Q sky130_fd_sc_hd__dfxtp_1
X_4459_ _5899_/S vssd1 vssd1 vccd1 vccd1 _5923_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7178_ _7178_/CLK _7178_/D vssd1 vssd1 vccd1 vccd1 _7178_/Q sky130_fd_sc_hd__dfxtp_1
X_6129_ _6129_/A _7649_/Q vssd1 vssd1 vccd1 vccd1 _6789_/A sky130_fd_sc_hd__xor2_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3072_ clkbuf_0__3072_/X vssd1 vssd1 vccd1 vccd1 _6246__398/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5681__239 _5681__239/A vssd1 vssd1 vccd1 vccd1 _7133_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _3738_/X _7587_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3831_/A sky130_fd_sc_hd__mux2_1
X_3761_ _3761_/A vssd1 vssd1 vccd1 vccd1 _7613_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3692_ _3707_/S vssd1 vssd1 vccd1 vccd1 _3701_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6480_ _6562_/A _6507_/B _6507_/C vssd1 vssd1 vccd1 vccd1 _6480_/Y sky130_fd_sc_hd__nand3b_1
X_5431_ _7177_/Q _7309_/Q _7495_/Q _7185_/Q _5252_/A _5397_/S vssd1 vssd1 vccd1 vccd1
+ _5431_/X sky130_fd_sc_hd__mux4_1
X_5362_ _7159_/Q _7151_/Q _5362_/S vssd1 vssd1 vccd1 vccd1 _5363_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7101_ _7525_/CLK _7101_/D vssd1 vssd1 vccd1 vccd1 _7101_/Q sky130_fd_sc_hd__dfxtp_1
X_4313_ _4313_/A vssd1 vssd1 vccd1 vccd1 _7371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5293_ _5293_/A _5292_/X vssd1 vssd1 vccd1 vccd1 _5293_/X sky130_fd_sc_hd__or2b_1
X_7032_ _7032_/A vssd1 vssd1 vccd1 vccd1 _7731_/D sky130_fd_sc_hd__clkbuf_1
X_4244_ _4243_/X _7398_/Q _4253_/S vssd1 vssd1 vccd1 vccd1 _4245_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3091_ _6333_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3091_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4175_ _4175_/A _4175_/B vssd1 vssd1 vccd1 vccd1 _4191_/S sky130_fd_sc_hd__or2_2
XFILLER_28_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6816_ _6816_/A _6816_/B vssd1 vssd1 vccd1 vccd1 _6817_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3959_ _3917_/X _7536_/Q _3963_/S vssd1 vssd1 vccd1 vccd1 _3960_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5629_ _7097_/Q _7196_/Q _5635_/S vssd1 vssd1 vccd1 vccd1 _5630_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6411__528 _6412__529/A vssd1 vssd1 vccd1 vccd1 _7470_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3289_ _6738_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3289_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2710_ clkbuf_0__2710_/X vssd1 vssd1 vccd1 vccd1 _5674__234/A sky130_fd_sc_hd__clkbuf_16
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3055_ clkbuf_0__3055_/X vssd1 vssd1 vccd1 vccd1 _6199__378/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6312__448 _6312__448/A vssd1 vssd1 vccd1 vccd1 _7390_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _7454_/Q _7446_/Q _7430_/Q _7422_/Q _5856_/X _5852_/X vssd1 vssd1 vccd1 vccd1
+ _5981_/B sky130_fd_sc_hd__mux4_1
XFILLER_18_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4931_ _4931_/A vssd1 vssd1 vccd1 vccd1 _7047_/D sky130_fd_sc_hd__clkbuf_1
X_4862_ _4843_/X _7114_/Q _4862_/S vssd1 vssd1 vccd1 vccd1 _4863_/A sky130_fd_sc_hd__mux2_1
X_7650_ _7655_/CLK _7650_/D vssd1 vssd1 vccd1 vccd1 _7650_/Q sky130_fd_sc_hd__dfxtp_1
X_3813_ _7669_/Q vssd1 vssd1 vccd1 vccd1 _3813_/X sky130_fd_sc_hd__buf_6
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6601_ _7512_/Q vssd1 vssd1 vccd1 vccd1 _6601_/Y sky130_fd_sc_hd__inv_2
X_7581_ _7581_/CLK _7581_/D vssd1 vssd1 vccd1 vccd1 _7581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4793_ _4793_/A vssd1 vssd1 vccd1 vccd1 _7142_/D sky130_fd_sc_hd__clkbuf_1
X_3744_ _3914_/A vssd1 vssd1 vccd1 vccd1 _3744_/X sky130_fd_sc_hd__buf_2
X_6532_ _6541_/B _6541_/C _6532_/C vssd1 vssd1 vccd1 vccd1 _6543_/B sky130_fd_sc_hd__and3_1
X_3675_ _3675_/A vssd1 vssd1 vccd1 vccd1 _7682_/D sky130_fd_sc_hd__clkbuf_1
X_6463_ _6463_/A _7513_/Q _6112_/A vssd1 vssd1 vccd1 vccd1 _6500_/A sky130_fd_sc_hd__or3b_1
Xoutput100 _5083_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[16] sky130_fd_sc_hd__buf_2
X_5414_ _7137_/Q _7060_/Q _7052_/Q _7273_/Q _5148_/A _5330_/S vssd1 vssd1 vccd1 vccd1
+ _5415_/B sky130_fd_sc_hd__mux4_1
Xoutput111 _5105_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput133 _4978_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput122 _4975_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[0] sky130_fd_sc_hd__buf_2
Xoutput155 _4967_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[1] sky130_fd_sc_hd__buf_2
Xoutput144 _4980_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput166 _5465_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput177 _5484_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[24] sky130_fd_sc_hd__buf_2
X_5345_ _7727_/Q vssd1 vssd1 vccd1 vccd1 _6149_/A sky130_fd_sc_hd__buf_2
Xoutput188 _5374_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[5] sky130_fd_sc_hd__buf_2
X_5276_ _7357_/Q _5339_/B _5469_/C vssd1 vssd1 vccd1 vccd1 _5276_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4227_ _4226_/X _7403_/Q _4227_/S vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__mux2_1
X_7015_ _6921_/A _6133_/A _7024_/S vssd1 vssd1 vccd1 vccd1 _7016_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3074_ _6254_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3074_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_68_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4158_ _4173_/S vssd1 vssd1 vccd1 vccd1 _4167_/S sky130_fd_sc_hd__buf_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4089_ _4089_/A vssd1 vssd1 vccd1 vccd1 _7458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5502__182 _5502__182/A vssd1 vssd1 vccd1 vccd1 _7038_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 caravel_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_2
Xinput24 caravel_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_2
Xinput35 caravel_wb_error_i vssd1 vssd1 vccd1 vccd1 _5492_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__3107_ clkbuf_0__3107_/X vssd1 vssd1 vccd1 vccd1 _6688_/A sky130_fd_sc_hd__clkbuf_16
Xinput46 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _5053_/A sky130_fd_sc_hd__buf_4
XFILLER_116_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput57 wbs_data_i[12] vssd1 vssd1 vccd1 vccd1 _5001_/A sky130_fd_sc_hd__buf_4
Xinput68 wbs_data_i[22] vssd1 vssd1 vccd1 vccd1 _5024_/A sky130_fd_sc_hd__buf_4
Xinput79 wbs_data_i[3] vssd1 vssd1 vccd1 vccd1 _3610_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5130_ _7350_/Q vssd1 vssd1 vccd1 vccd1 _5205_/A sky130_fd_sc_hd__clkinv_2
X_5061_ _5061_/A vssd1 vssd1 vccd1 vccd1 _5061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4012_ _4012_/A vssd1 vssd1 vccd1 vccd1 _7492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2967_ clkbuf_0__2967_/X vssd1 vssd1 vccd1 vccd1 _6173__357/A sky130_fd_sc_hd__clkbuf_16
XFILLER_53_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5963_ _7397_/Q _7239_/Q _7555_/Q _7461_/Q _5925_/A _4468_/A vssd1 vssd1 vccd1 vccd1
+ _5964_/B sky130_fd_sc_hd__mux4_1
XFILLER_92_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7702_ _7702_/CLK _7702_/D vssd1 vssd1 vccd1 vccd1 _7702_/Q sky130_fd_sc_hd__dfxtp_1
X_4914_ _4840_/X _7054_/Q _4916_/S vssd1 vssd1 vccd1 vccd1 _4915_/A sky130_fd_sc_hd__mux2_1
X_5894_ _7536_/Q _7677_/Q _7693_/Q _7279_/Q _5884_/A _4462_/A vssd1 vssd1 vccd1 vccd1
+ _5894_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7633_ _7633_/CLK _7633_/D vssd1 vssd1 vccd1 vccd1 _7633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2712_ _5676_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2712_/X sky130_fd_sc_hd__clkbuf_16
X_4845_ _4845_/A vssd1 vssd1 vccd1 vccd1 _7122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7564_ _7564_/CLK _7564_/D vssd1 vssd1 vccd1 vccd1 _7564_/Q sky130_fd_sc_hd__dfxtp_2
X_4776_ _7149_/Q _4334_/X _4782_/S vssd1 vssd1 vccd1 vccd1 _4777_/A sky130_fd_sc_hd__mux2_1
X_3727_ _3727_/A vssd1 vssd1 vccd1 vccd1 _7623_/D sky130_fd_sc_hd__clkbuf_1
X_6515_ _6515_/A _6515_/B _7514_/Q vssd1 vssd1 vccd1 vccd1 _6515_/X sky130_fd_sc_hd__or3b_1
X_7495_ _7495_/CLK _7495_/D vssd1 vssd1 vccd1 vccd1 _7495_/Q sky130_fd_sc_hd__dfxtp_1
X_3658_ _3658_/A vssd1 vssd1 vccd1 vccd1 _7686_/D sky130_fd_sc_hd__clkbuf_1
X_6446_ _6446_/A _6446_/B _6093_/Y vssd1 vssd1 vccd1 vccd1 _6448_/B sky130_fd_sc_hd__or3b_1
XFILLER_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3589_ _7704_/Q _3588_/X _3595_/S vssd1 vssd1 vccd1 vccd1 _3590_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5328_ _5264_/X _5327_/X _4368_/A vssd1 vssd1 vccd1 vccd1 _5328_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5259_ _5259_/A vssd1 vssd1 vccd1 vccd1 _5259_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_0__3057_ _6207_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3057_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6051__331 _6052__332/A vssd1 vssd1 vccd1 vccd1 _7257_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _4246_/X _7247_/Q _4634_/S vssd1 vssd1 vccd1 vccd1 _4631_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4561_ _4561_/A _4561_/B _4301_/A vssd1 vssd1 vccd1 vccd1 _4918_/B sky130_fd_sc_hd__or3b_4
XFILLER_116_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7280_ _7280_/CLK _7280_/D vssd1 vssd1 vccd1 vccd1 _7280_/Q sky130_fd_sc_hd__dfxtp_1
X_4492_ _4217_/X _7308_/Q _4498_/S vssd1 vssd1 vccd1 vccd1 _4493_/A sky130_fd_sc_hd__mux2_1
X_3512_ _5185_/B _3501_/X _5586_/C _3510_/X _5587_/B vssd1 vssd1 vccd1 vccd1 _3513_/A
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6231_ _7666_/Q _6231_/B vssd1 vssd1 vccd1 vccd1 _6232_/A sky130_fd_sc_hd__and2_1
XFILLER_103_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3097_ clkbuf_0__3097_/X vssd1 vssd1 vccd1 vccd1 _6369__494/A sky130_fd_sc_hd__clkbuf_16
X_6162_ _7720_/Q _7651_/Q vssd1 vssd1 vccd1 vccd1 _6791_/C sky130_fd_sc_hd__xor2_1
XFILLER_97_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _7083_/Q _7084_/Q vssd1 vssd1 vccd1 vccd1 _5232_/A sky130_fd_sc_hd__or2_2
X_5702__256 _5702__256/A vssd1 vssd1 vccd1 vccd1 _7150_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _7723_/Q _6129_/A vssd1 vssd1 vccd1 vccd1 _6093_/Y sky130_fd_sc_hd__nor2_1
X_5044_ _5044_/A _5046_/B vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__and2_1
XFILLER_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6995_ _7031_/A _6995_/B vssd1 vssd1 vccd1 vccd1 _6996_/A sky130_fd_sc_hd__or2_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5946_ _7626_/Q _7618_/Q _7602_/Q _7594_/Q _5870_/X _5925_/X vssd1 vssd1 vccd1 vccd1
+ _5947_/B sky130_fd_sc_hd__mux4_2
XFILLER_53_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5877_ _7314_/Q vssd1 vssd1 vccd1 vccd1 _5882_/A sky130_fd_sc_hd__clkbuf_2
X_7616_ _7616_/CLK _7616_/D vssd1 vssd1 vccd1 vccd1 _7616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4828_ _7326_/Q vssd1 vssd1 vccd1 vccd1 _4828_/X sky130_fd_sc_hd__buf_2
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7547_ _7547_/CLK _7547_/D vssd1 vssd1 vccd1 vccd1 _7547_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__2626_ _5497_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2626_/X sky130_fd_sc_hd__clkbuf_16
X_4759_ _4759_/A vssd1 vssd1 vccd1 vccd1 _7158_/D sky130_fd_sc_hd__clkbuf_1
X_7478_ _7478_/CLK _7478_/D vssd1 vssd1 vccd1 vccd1 _7478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3109_ _6421_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3109_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_76_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _3652_/X _7521_/Q _3994_/S vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6780_ _6878_/A _6878_/B _6878_/D vssd1 vssd1 vccd1 vccd1 _6780_/Y sky130_fd_sc_hd__nor3_1
XFILLER_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5800_ _7209_/Q _5044_/A _5800_/S vssd1 vssd1 vccd1 vccd1 _5801_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2666_ clkbuf_0__2666_/X vssd1 vssd1 vccd1 vccd1 _5650__214/A sky130_fd_sc_hd__clkbuf_16
X_5731_ _5731_/A vssd1 vssd1 vccd1 vccd1 _5731_/X sky130_fd_sc_hd__buf_1
X_4613_ _4613_/A vssd1 vssd1 vccd1 vccd1 _7255_/D sky130_fd_sc_hd__clkbuf_1
X_7401_ _7401_/CLK _7401_/D vssd1 vssd1 vccd1 vccd1 _7401_/Q sky130_fd_sc_hd__dfxtp_2
X_5593_ _5637_/A vssd1 vssd1 vccd1 vccd1 _5602_/S sky130_fd_sc_hd__buf_2
X_4544_ _7284_/Q _3899_/A _4552_/S vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__mux2_1
X_7332_ _7332_/CLK _7332_/D vssd1 vssd1 vccd1 vccd1 _7332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7263_ _7263_/CLK _7263_/D vssd1 vssd1 vccd1 vccd1 _7263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4475_ _4475_/A vssd1 vssd1 vccd1 vccd1 _7313_/D sky130_fd_sc_hd__clkbuf_1
X_6214_ _6214_/A vssd1 vssd1 vccd1 vccd1 _6214_/X sky130_fd_sc_hd__buf_1
X_7194_ _7727_/CLK _7194_/D vssd1 vssd1 vccd1 vccd1 _7194_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6145_ _6144_/Y _7640_/Q _6143_/B vssd1 vssd1 vccd1 vccd1 _6788_/A sky130_fd_sc_hd__o21a_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_15 _5495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6076_ _7276_/Q _5766_/A _6076_/S vssd1 vssd1 vccd1 vccd1 _6077_/A sky130_fd_sc_hd__mux2_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _5027_/A _5035_/B vssd1 vssd1 vccd1 vccd1 _5028_/A sky130_fd_sc_hd__and2_1
XINSDIODE2_59 _3914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_26 _7557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_48 _3549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_37 _5049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6978_ _5010_/A _7716_/Q _6978_/S vssd1 vssd1 vccd1 vccd1 _6979_/B sky130_fd_sc_hd__mux2_1
X_5929_ _5929_/A vssd1 vssd1 vccd1 vccd1 _5929_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6742__173 _6743__174/A vssd1 vssd1 vccd1 vccd1 _7617_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__3286_ clkbuf_0__3286_/X vssd1 vssd1 vccd1 vccd1 _6724__158/A sky130_fd_sc_hd__clkbuf_16
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4260_ _4260_/A vssd1 vssd1 vccd1 vccd1 _7393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4191_ _4118_/X _7416_/Q _4191_/S vssd1 vssd1 vccd1 vccd1 _4192_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__2960_ _6056_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2960_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6901_ _7664_/Q _6905_/B vssd1 vssd1 vccd1 vccd1 _6901_/X sky130_fd_sc_hd__or2_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6832_ _6832_/A vssd1 vssd1 vccd1 vccd1 _7645_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2718_ clkbuf_0__2718_/X vssd1 vssd1 vccd1 vccd1 _5712__264/A sky130_fd_sc_hd__clkbuf_16
X_3975_ _3656_/X _7529_/Q _3975_/S vssd1 vssd1 vccd1 vccd1 _3976_/A sky130_fd_sc_hd__mux2_1
X_6763_ _6763_/A vssd1 vssd1 vccd1 vccd1 _6763_/X sky130_fd_sc_hd__buf_1
X_6064__341 _6065__342/A vssd1 vssd1 vccd1 vccd1 _7267_/CLK sky130_fd_sc_hd__inv_2
X_5645_ _5645_/A _5645_/B vssd1 vssd1 vccd1 vccd1 _5645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7315_ _7315_/CLK _7315_/D vssd1 vssd1 vccd1 vccd1 _7315_/Q sky130_fd_sc_hd__dfxtp_1
X_4527_ _4527_/A vssd1 vssd1 vccd1 vccd1 _7293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7246_ _7246_/CLK _7246_/D vssd1 vssd1 vccd1 vccd1 _7246_/Q sky130_fd_sc_hd__dfxtp_1
X_4458_ _5869_/A vssd1 vssd1 vccd1 vccd1 _5899_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_6685__127 _6685__127/A vssd1 vssd1 vccd1 vccd1 _7571_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7177_ _7177_/CLK _7177_/D vssd1 vssd1 vccd1 vccd1 _7177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6128_ _6128_/A vssd1 vssd1 vccd1 vccd1 _6777_/A sky130_fd_sc_hd__clkbuf_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4389_ _4384_/A _4391_/B _4388_/Y vssd1 vssd1 vccd1 vccd1 _7350_/D sky130_fd_sc_hd__o21a_1
XFILLER_105_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5715__266 _5716__267/A vssd1 vssd1 vccd1 vccd1 _7160_/CLK sky130_fd_sc_hd__inv_2
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3760_ _3633_/X _7613_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3761_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__3269_ clkbuf_0__3269_/X vssd1 vssd1 vccd1 vccd1 _6637__88/A sky130_fd_sc_hd__clkbuf_16
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3691_ _4283_/A _4175_/A vssd1 vssd1 vccd1 vccd1 _3707_/S sky130_fd_sc_hd__or2_2
X_5430_ _5252_/X _5429_/X _5213_/A vssd1 vssd1 vccd1 vccd1 _5430_/X sky130_fd_sc_hd__a21o_1
X_5361_ _5363_/A _5358_/Y _5360_/Y _5415_/A vssd1 vssd1 vccd1 vccd1 _5361_/X sky130_fd_sc_hd__o211a_1
X_5292_ _7520_/Q _7141_/Q _5299_/A vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__mux2_1
X_7100_ _7727_/CLK _7100_/D vssd1 vssd1 vccd1 vccd1 _7100_/Q sky130_fd_sc_hd__dfxtp_1
X_4312_ _4226_/X _7371_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4243_ _7673_/Q vssd1 vssd1 vccd1 vccd1 _4243_/X sky130_fd_sc_hd__clkbuf_4
X_7031_ _7031_/A _7031_/B vssd1 vssd1 vccd1 vccd1 _7032_/A sky130_fd_sc_hd__or2_1
XFILLER_101_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6749__179 _6749__179/A vssd1 vssd1 vccd1 vccd1 _7623_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3090_ _6327_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3090_/X sky130_fd_sc_hd__clkbuf_16
X_4174_ _4174_/A vssd1 vssd1 vccd1 vccd1 _7424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6636__87 _6638__89/A vssd1 vssd1 vccd1 vccd1 _7531_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6815_ _6816_/A _6816_/B vssd1 vssd1 vccd1 vccd1 _6821_/B sky130_fd_sc_hd__nor2_1
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6691__131 _6691__131/A vssd1 vssd1 vccd1 vccd1 _7575_/CLK sky130_fd_sc_hd__inv_2
X_3958_ _3958_/A vssd1 vssd1 vccd1 vccd1 _7537_/D sky130_fd_sc_hd__clkbuf_1
X_3889_ _7562_/Q _3591_/X _3891_/S vssd1 vssd1 vccd1 vccd1 _3890_/A sky130_fd_sc_hd__mux2_1
X_5628_ _5628_/A vssd1 vssd1 vccd1 vccd1 _7096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5559_ _5642_/A vssd1 vssd1 vccd1 vccd1 _5645_/A sky130_fd_sc_hd__inv_2
XFILLER_105_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7229_ _7229_/CLK _7229_/D vssd1 vssd1 vccd1 vccd1 _7229_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3288_ _6732_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3288_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_100_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6379__502 _6379__502/A vssd1 vssd1 vccd1 vccd1 _7444_/CLK sky130_fd_sc_hd__inv_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__3054_ clkbuf_0__3054_/X vssd1 vssd1 vccd1 vccd1 _6194__374/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6015__302 _6015__302/A vssd1 vssd1 vccd1 vccd1 _7228_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4930_ _7047_/Q _4578_/A _4934_/S vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4861_ _4861_/A vssd1 vssd1 vccd1 vccd1 _7115_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3812_ _3812_/A vssd1 vssd1 vccd1 vccd1 _7593_/D sky130_fd_sc_hd__clkbuf_1
X_6600_ _6600_/A vssd1 vssd1 vccd1 vccd1 _7511_/D sky130_fd_sc_hd__clkbuf_1
X_7580_ _7580_/CLK _7580_/D vssd1 vssd1 vccd1 vccd1 _7580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4792_ _7142_/Q _4572_/A _4794_/S vssd1 vssd1 vccd1 vccd1 _4793_/A sky130_fd_sc_hd__mux2_1
X_3743_ _3743_/A vssd1 vssd1 vccd1 vccd1 _7618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6531_ _6529_/Y _6526_/X _6530_/X _5991_/X vssd1 vssd1 vccd1 vccd1 _7499_/D sky130_fd_sc_hd__o211a_1
X_3674_ _3469_/X _7682_/Q _3682_/S vssd1 vssd1 vccd1 vccd1 _3675_/A sky130_fd_sc_hd__mux2_1
X_6462_ _6462_/A _6462_/B vssd1 vssd1 vccd1 vccd1 _6503_/B sky130_fd_sc_hd__xnor2_2
Xoutput101 _5085_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[17] sky130_fd_sc_hd__buf_2
X_5413_ _5413_/A _5413_/B vssd1 vssd1 vccd1 vccd1 _5413_/X sky130_fd_sc_hd__or2_1
Xoutput112 _5107_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[27] sky130_fd_sc_hd__buf_2
Xoutput134 _5021_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[20] sky130_fd_sc_hd__buf_2
Xoutput123 _4998_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[10] sky130_fd_sc_hd__buf_2
X_5344_ _5458_/A _7066_/Q _5376_/A input30/X vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__a22o_1
Xoutput145 _5043_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[30] sky130_fd_sc_hd__buf_2
Xoutput156 _4971_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[2] sky130_fd_sc_hd__buf_2
Xoutput167 _5468_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput189 _5411_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[6] sky130_fd_sc_hd__buf_2
Xoutput178 _5485_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[25] sky130_fd_sc_hd__buf_2
X_5275_ _5337_/A _5255_/X _5274_/X _5308_/A vssd1 vssd1 vccd1 vccd1 _5275_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4226_ _4575_/A vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__clkbuf_4
X_7014_ _7014_/A vssd1 vssd1 vccd1 vccd1 _7725_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3073_ _6248_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3073_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4157_ _4642_/A _4175_/B vssd1 vssd1 vccd1 vccd1 _4173_/S sky130_fd_sc_hd__or2_2
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4088_ _7458_/Q _3813_/X _4092_/S vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__mux2_1
X_6624__79 _6624__79/A vssd1 vssd1 vccd1 vccd1 _7522_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6374__498 _6375__499/A vssd1 vssd1 vccd1 vccd1 _7440_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6698__137 _6698__137/A vssd1 vssd1 vccd1 vccd1 _7581_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput25 caravel_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_4
Xinput14 caravel_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__3106_ clkbuf_0__3106_/X vssd1 vssd1 vccd1 vccd1 _6418__534/A sky130_fd_sc_hd__clkbuf_16
Xinput36 wb_rst_i vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__buf_4
Xinput69 wbs_data_i[23] vssd1 vssd1 vccd1 vccd1 _5027_/A sky130_fd_sc_hd__buf_4
Xinput58 wbs_data_i[13] vssd1 vssd1 vccd1 vccd1 _5004_/A sky130_fd_sc_hd__buf_4
XFILLER_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5060_ _5060_/A _5068_/B vssd1 vssd1 vccd1 vccd1 _5061_/A sky130_fd_sc_hd__and2_1
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4011_ _7492_/Q _3591_/X _4013_/S vssd1 vssd1 vccd1 vccd1 _4012_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2966_ clkbuf_0__2966_/X vssd1 vssd1 vccd1 vccd1 _6085__354/A sky130_fd_sc_hd__clkbuf_16
XFILLER_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5962_ _6001_/A _5962_/B vssd1 vssd1 vccd1 vccd1 _5962_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7701_ _7701_/CLK _7701_/D vssd1 vssd1 vccd1 vccd1 _7701_/Q sky130_fd_sc_hd__dfxtp_1
X_4913_ _4913_/A vssd1 vssd1 vccd1 vccd1 _7055_/D sky130_fd_sc_hd__clkbuf_1
X_5893_ _4473_/A _5886_/Y _5888_/Y _5890_/Y _5892_/Y vssd1 vssd1 vccd1 vccd1 _5893_/X
+ sky130_fd_sc_hd__o32a_1
X_7632_ _7632_/CLK _7632_/D vssd1 vssd1 vccd1 vccd1 _7632_/Q sky130_fd_sc_hd__dfxtp_1
X_4844_ _4843_/X _7122_/Q _4844_/S vssd1 vssd1 vccd1 vccd1 _4845_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2711_ _5675_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2711_/X sky130_fd_sc_hd__clkbuf_16
X_7563_ _7563_/CLK _7563_/D vssd1 vssd1 vccd1 vccd1 _7563_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4775_ _4775_/A vssd1 vssd1 vccd1 vccd1 _7150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3726_ _3542_/X _7623_/Q _3728_/S vssd1 vssd1 vccd1 vccd1 _3727_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6514_ _7515_/Q vssd1 vssd1 vccd1 vccd1 _6515_/B sky130_fd_sc_hd__inv_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7494_ _7494_/CLK _7494_/D vssd1 vssd1 vccd1 vccd1 _7494_/Q sky130_fd_sc_hd__dfxtp_1
X_3657_ _3656_/X _7686_/Q _3657_/S vssd1 vssd1 vccd1 vccd1 _3658_/A sky130_fd_sc_hd__mux2_1
X_6445_ _7509_/Q _6445_/B vssd1 vssd1 vccd1 vccd1 _6504_/D sky130_fd_sc_hd__xnor2_1
X_6376_ _6382_/A vssd1 vssd1 vccd1 vccd1 _6376_/X sky130_fd_sc_hd__buf_1
X_3588_ _7326_/Q vssd1 vssd1 vccd1 vccd1 _3588_/X sky130_fd_sc_hd__buf_4
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5327_ _7372_/Q _7343_/Q _7335_/Q _7298_/Q _5325_/S _5210_/A vssd1 vssd1 vccd1 vccd1
+ _5327_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5258_ _7116_/Q _7164_/Q _5421_/S vssd1 vssd1 vccd1 vccd1 _5259_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3056_ _6201_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3056_/X sky130_fd_sc_hd__clkbuf_16
X_4209_ _4118_/X _7408_/Q _4209_/S vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5189_ _5162_/X _5181_/X _5184_/Y _5339_/B vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__a31o_1
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6754__7 _6754__7/A vssd1 vssd1 vccd1 vccd1 _7626_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6706__144 _6706__144/A vssd1 vssd1 vccd1 vccd1 _7588_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4560_/A vssd1 vssd1 vccd1 vccd1 _4560_/X sky130_fd_sc_hd__buf_2
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4491_ _4491_/A vssd1 vssd1 vccd1 vccd1 _7309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3511_ _3511_/A _6910_/B vssd1 vssd1 vccd1 vccd1 _5587_/B sky130_fd_sc_hd__or2b_4
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6230_ _6230_/A vssd1 vssd1 vccd1 vccd1 _7327_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__3096_ clkbuf_0__3096_/X vssd1 vssd1 vccd1 vccd1 _6360__486/A sky130_fd_sc_hd__clkbuf_16
XFILLER_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6462_/B _6161_/B vssd1 vssd1 vccd1 vccd1 _6774_/B sky130_fd_sc_hd__xnor2_1
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5112_/A vssd1 vssd1 vccd1 vccd1 _5112_/X sky130_fd_sc_hd__clkbuf_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _7727_/Q _7726_/Q _7725_/Q _7724_/Q vssd1 vssd1 vccd1 vccd1 _6127_/C sky130_fd_sc_hd__or4_2
X_5043_ _5043_/A vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__clkbuf_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6994_ _5001_/A _7720_/Q _7007_/S vssd1 vssd1 vccd1 vccd1 _6995_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6028__312 _6030__314/A vssd1 vssd1 vccd1 vccd1 _7238_/CLK sky130_fd_sc_hd__inv_2
X_5945_ _6003_/A _5945_/B vssd1 vssd1 vccd1 vccd1 _5945_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6325__459 _6325__459/A vssd1 vssd1 vccd1 vccd1 _7401_/CLK sky130_fd_sc_hd__inv_2
X_5876_ _6001_/A _5873_/X _5875_/X _5917_/A vssd1 vssd1 vccd1 vccd1 _5876_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7615_ _7615_/CLK _7615_/D vssd1 vssd1 vccd1 vccd1 _7615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4827_ _4827_/A vssd1 vssd1 vccd1 vccd1 _7128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7546_ _7546_/CLK _7546_/D vssd1 vssd1 vccd1 vccd1 _7546_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__2625_ _5496_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2625_/X sky130_fd_sc_hd__clkbuf_16
X_4758_ _4572_/X _7158_/Q _4760_/S vssd1 vssd1 vccd1 vccd1 _4759_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4689_ _4689_/A vssd1 vssd1 vccd1 vccd1 _7213_/D sky130_fd_sc_hd__clkbuf_1
X_7477_ _7477_/CLK _7477_/D vssd1 vssd1 vccd1 vccd1 _7477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3709_ _7318_/Q vssd1 vssd1 vccd1 vccd1 _4587_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3108_ _6420_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3108_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_17_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3991_ _3991_/A vssd1 vssd1 vccd1 vccd1 _7522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__2665_ clkbuf_0__2665_/X vssd1 vssd1 vccd1 vccd1 _5663_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7400_ _7400_/CLK _7400_/D vssd1 vssd1 vccd1 vccd1 _7400_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4612_ _7255_/Q _3908_/A _4616_/S vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__mux2_1
X_5592_ _5535_/B _5645_/B _5643_/B _5592_/D vssd1 vssd1 vccd1 vccd1 _5637_/A sky130_fd_sc_hd__and4b_4
X_4543_ _4558_/S vssd1 vssd1 vccd1 vccd1 _4552_/S sky130_fd_sc_hd__clkbuf_2
X_7331_ _7331_/CLK _7331_/D vssd1 vssd1 vccd1 vccd1 _7331_/Q sky130_fd_sc_hd__dfxtp_1
X_7262_ _7262_/CLK _7262_/D vssd1 vssd1 vccd1 vccd1 _7262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4474_ _4486_/C _4474_/B _4474_/C vssd1 vssd1 vccd1 vccd1 _4475_/A sky130_fd_sc_hd__and3_1
X_7193_ _7722_/CLK _7193_/D vssd1 vssd1 vccd1 vccd1 _7193_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_97_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6144_ _6487_/A vssd1 vssd1 vccd1 vccd1 _6144_/Y sky130_fd_sc_hd__inv_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_16 _5873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6331__463 _6331__463/A vssd1 vssd1 vccd1 vccd1 _7405_/CLK sky130_fd_sc_hd__inv_2
X_6075_ _6075_/A vssd1 vssd1 vccd1 vccd1 _7275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_38 _5053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5026_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5035_/B sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_27 _7041_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6972__4 _6972__4/A vssd1 vssd1 vccd1 vccd1 _7714_/CLK sky130_fd_sc_hd__inv_2
XINSDIODE2_49 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6977_ _6977_/A vssd1 vssd1 vccd1 vccd1 _7715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5928_ _7411_/Q _7379_/Q _7710_/Q _7633_/Q _5819_/X _4484_/X vssd1 vssd1 vccd1 vccd1
+ _5928_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5859_ _6005_/A _5858_/X _3485_/Y vssd1 vssd1 vccd1 vccd1 _5859_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7529_ _7529_/CLK _7529_/D vssd1 vssd1 vccd1 vccd1 _7529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__3285_ clkbuf_0__3285_/X vssd1 vssd1 vccd1 vccd1 _6744_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4190_ _4190_/A vssd1 vssd1 vccd1 vccd1 _7417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6900_ _7663_/Q _6893_/B _6899_/X _6886_/X vssd1 vssd1 vccd1 vccd1 _7663_/D sky130_fd_sc_hd__o211a_1
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6831_ _6835_/B _6831_/B _6872_/B vssd1 vssd1 vccd1 vccd1 _6832_/A sky130_fd_sc_hd__and3b_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2717_ clkbuf_0__2717_/X vssd1 vssd1 vccd1 vccd1 _5725_/A sky130_fd_sc_hd__clkbuf_16
X_3974_ _3974_/A vssd1 vssd1 vccd1 vccd1 _7530_/D sky130_fd_sc_hd__clkbuf_1
X_6209__385 _6210__386/A vssd1 vssd1 vccd1 vccd1 _7315_/CLK sky130_fd_sc_hd__inv_2
X_5713_ _5725_/A vssd1 vssd1 vccd1 vccd1 _5713_/X sky130_fd_sc_hd__buf_1
X_5644_ _3511_/A _6910_/B _5590_/A _5642_/Y _5647_/B vssd1 vssd1 vccd1 vccd1 _7103_/D
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_117_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7314_ _7314_/CLK _7314_/D vssd1 vssd1 vccd1 vccd1 _7314_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_4_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5496_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4526_ _4211_/X _7293_/Q _4534_/S vssd1 vssd1 vccd1 vccd1 _4527_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7245_ _7245_/CLK _7245_/D vssd1 vssd1 vccd1 vccd1 _7245_/Q sky130_fd_sc_hd__dfxtp_1
X_4457_ _7312_/Q vssd1 vssd1 vccd1 vccd1 _5869_/A sky130_fd_sc_hd__buf_2
X_6175__359 _6175__359/A vssd1 vssd1 vccd1 vccd1 _7289_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7176_ _7176_/CLK _7176_/D vssd1 vssd1 vccd1 vccd1 _7176_/Q sky130_fd_sc_hd__dfxtp_1
X_6127_ _7723_/Q _6127_/B _6127_/C vssd1 vssd1 vccd1 vccd1 _6128_/A sky130_fd_sc_hd__or3_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4388_ _6274_/A _4388_/B vssd1 vssd1 vccd1 vccd1 _4388_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5009_ _5009_/A vssd1 vssd1 vccd1 vccd1 _5009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6338__469 _6338__469/A vssd1 vssd1 vccd1 vccd1 _7411_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3268_ clkbuf_0__3268_/X vssd1 vssd1 vccd1 vccd1 _6628__81/A sky130_fd_sc_hd__clkbuf_16
XFILLER_9_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3690_ _3484_/A _3796_/C _4606_/A vssd1 vssd1 vccd1 vccd1 _4175_/A sky130_fd_sc_hd__nand3b_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5360_ _5360_/A _5360_/B vssd1 vssd1 vccd1 vccd1 _5360_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5291_ _5291_/A _5291_/B vssd1 vssd1 vccd1 vccd1 _5291_/Y sky130_fd_sc_hd__nand2_1
X_4311_ _4311_/A vssd1 vssd1 vccd1 vccd1 _7372_/D sky130_fd_sc_hd__clkbuf_1
X_4242_ _4242_/A vssd1 vssd1 vccd1 vccd1 _7399_/D sky130_fd_sc_hd__clkbuf_1
X_7030_ _6911_/A _5235_/X _7033_/S vssd1 vssd1 vccd1 vccd1 _7031_/B sky130_fd_sc_hd__mux2_1
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4173_ _4118_/X _7424_/Q _4173_/S vssd1 vssd1 vccd1 vccd1 _4174_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6814_ _6814_/A vssd1 vssd1 vccd1 vccd1 _7641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3957_ _3914_/X _7537_/Q _3957_/S vssd1 vssd1 vccd1 vccd1 _3958_/A sky130_fd_sc_hd__mux2_1
X_6181__363 _6182__364/A vssd1 vssd1 vccd1 vccd1 _7293_/CLK sky130_fd_sc_hd__inv_2
X_6676_ _6682_/A vssd1 vssd1 vccd1 vccd1 _6676_/X sky130_fd_sc_hd__buf_1
X_3888_ _3888_/A vssd1 vssd1 vccd1 vccd1 _7563_/D sky130_fd_sc_hd__clkbuf_1
X_5627_ _7096_/Q _7195_/Q _5635_/S vssd1 vssd1 vccd1 vccd1 _5628_/A sky130_fd_sc_hd__mux2_1
X_5558_ _7070_/Q _7069_/Q _5642_/A _5557_/X vssd1 vssd1 vccd1 vccd1 _7069_/D sky130_fd_sc_hd__o31a_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4509_ _4509_/A vssd1 vssd1 vccd1 vccd1 _7301_/D sky130_fd_sc_hd__clkbuf_1
X_7228_ _7228_/CLK _7228_/D vssd1 vssd1 vccd1 vccd1 _7228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5489_ _5375_/X _7207_/Q input24/X _5376_/X vssd1 vssd1 vccd1 vccd1 _5489_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3287_ _6726_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3287_/X sky130_fd_sc_hd__clkbuf_16
X_5721__271 _5723__273/A vssd1 vssd1 vccd1 vccd1 _7165_/CLK sky130_fd_sc_hd__inv_2
X_7159_ _7159_/CLK _7159_/D vssd1 vssd1 vccd1 vccd1 _7159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6700__139 _6700__139/A vssd1 vssd1 vccd1 vccd1 _7583_/CLK sky130_fd_sc_hd__inv_2
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3053_ clkbuf_0__3053_/X vssd1 vssd1 vccd1 vccd1 _6186__367/A sky130_fd_sc_hd__clkbuf_16
XFILLER_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5577__208 _5578__209/A vssd1 vssd1 vccd1 vccd1 _7076_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6641__91 _6644__94/A vssd1 vssd1 vccd1 vccd1 _7535_/CLK sky130_fd_sc_hd__inv_2
X_4860_ _4840_/X _7115_/Q _4862_/S vssd1 vssd1 vccd1 vccd1 _4861_/A sky130_fd_sc_hd__mux2_1
X_3811_ _7593_/Q _3810_/X _3811_/S vssd1 vssd1 vccd1 vccd1 _3812_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4791_ _4791_/A vssd1 vssd1 vccd1 vccd1 _7143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6530_ _6532_/C _6566_/A _6541_/C vssd1 vssd1 vccd1 vccd1 _6530_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3742_ _3741_/X _7618_/Q _3745_/S vssd1 vssd1 vccd1 vccd1 _3743_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3673_ _3688_/S vssd1 vssd1 vccd1 vccd1 _3682_/S sky130_fd_sc_hd__buf_2
X_5664__225 _5668__229/A vssd1 vssd1 vccd1 vccd1 _7119_/CLK sky130_fd_sc_hd__inv_2
X_6461_ _7510_/Q vssd1 vssd1 vccd1 vccd1 _6594_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5412_ _7549_/Q _7439_/Q _7407_/Q _7391_/Q _5285_/S _5210_/A vssd1 vssd1 vccd1 vccd1
+ _5413_/B sky130_fd_sc_hd__mux4_2
Xoutput102 _5087_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput113 _5052_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[2] sky130_fd_sc_hd__buf_2
Xoutput124 _5000_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[11] sky130_fd_sc_hd__buf_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5343_ _5343_/A _5343_/B vssd1 vssd1 vccd1 vccd1 _5343_/Y sky130_fd_sc_hd__nand2_1
Xoutput146 _5045_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[31] sky130_fd_sc_hd__buf_2
Xoutput135 _5023_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[21] sky130_fd_sc_hd__buf_2
Xoutput157 _4973_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[3] sky130_fd_sc_hd__buf_2
Xoutput168 _5471_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_102_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput179 _5486_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[26] sky130_fd_sc_hd__buf_2
X_5274_ _5158_/X _5257_/Y _5263_/X _5273_/X _5161_/A vssd1 vssd1 vccd1 vccd1 _5274_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4225_ _4225_/A vssd1 vssd1 vccd1 vccd1 _7404_/D sky130_fd_sc_hd__clkbuf_1
X_7013_ _7003_/X _7013_/B vssd1 vssd1 vccd1 vccd1 _7014_/A sky130_fd_sc_hd__and2b_1
Xclkbuf_0__3072_ _6242_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3072_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_110_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4156_ _4156_/A vssd1 vssd1 vccd1 vccd1 _7432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _4087_/A vssd1 vssd1 vccd1 vccd1 _7459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4989_ _4989_/A vssd1 vssd1 vccd1 vccd1 _4989_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6188__369 _6188__369/A vssd1 vssd1 vccd1 vccd1 _7299_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3105_ clkbuf_0__3105_/X vssd1 vssd1 vccd1 vccd1 _6412__529/A sky130_fd_sc_hd__clkbuf_16
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput26 caravel_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_2
Xinput15 caravel_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_2
Xinput37 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__buf_4
XFILLER_116_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput48 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _5057_/A sky130_fd_sc_hd__buf_4
Xinput59 wbs_data_i[14] vssd1 vssd1 vccd1 vccd1 _5006_/A sky130_fd_sc_hd__buf_4
X_5728__277 _5728__277/A vssd1 vssd1 vccd1 vccd1 _7171_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4010_ _4010_/A vssd1 vssd1 vccd1 vccd1 _7493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5961_ _7453_/Q _7445_/Q _7429_/Q _7421_/Q _5856_/X _5852_/X vssd1 vssd1 vccd1 vccd1
+ _5962_/B sky130_fd_sc_hd__mux4_1
X_7700_ _7700_/CLK _7700_/D vssd1 vssd1 vccd1 vccd1 _7700_/Q sky130_fd_sc_hd__dfxtp_1
X_4912_ _4837_/X _7055_/Q _4916_/S vssd1 vssd1 vccd1 vccd1 _4913_/A sky130_fd_sc_hd__mux2_1
X_7631_ _7631_/CLK _7631_/D vssd1 vssd1 vccd1 vccd1 _7631_/Q sky130_fd_sc_hd__dfxtp_1
X_5892_ _5888_/A _5891_/X _4473_/A vssd1 vssd1 vccd1 vccd1 _5892_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2710_ _5669_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2710_/X sky130_fd_sc_hd__clkbuf_16
X_4843_ _7321_/Q vssd1 vssd1 vccd1 vccd1 _4843_/X sky130_fd_sc_hd__buf_2
X_7562_ _7562_/CLK _7562_/D vssd1 vssd1 vccd1 vccd1 _7562_/Q sky130_fd_sc_hd__dfxtp_2
X_4774_ _7150_/Q _4331_/X _4774_/S vssd1 vssd1 vccd1 vccd1 _4775_/A sky130_fd_sc_hd__mux2_1
X_3725_ _3725_/A vssd1 vssd1 vccd1 vccd1 _7624_/D sky130_fd_sc_hd__clkbuf_1
X_7493_ _7493_/CLK _7493_/D vssd1 vssd1 vccd1 vccd1 _7493_/Q sky130_fd_sc_hd__dfxtp_1
X_6513_ _7516_/Q vssd1 vssd1 vccd1 vccd1 _6515_/A sky130_fd_sc_hd__inv_2
X_6444_ _7720_/Q _6163_/A _6462_/B vssd1 vssd1 vccd1 vccd1 _6445_/B sky130_fd_sc_hd__a21oi_1
X_3656_ _4575_/A vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__buf_2
X_3587_ _3587_/A vssd1 vssd1 vccd1 vccd1 _7705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5326_ _5360_/A _5325_/X vssd1 vssd1 vccd1 vccd1 _5326_/X sky130_fd_sc_hd__or2b_1
XFILLER_102_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5525__195 _5528__198/A vssd1 vssd1 vccd1 vccd1 _7052_/CLK sky130_fd_sc_hd__inv_2
X_5257_ _5257_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5257_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4208_ _4208_/A vssd1 vssd1 vccd1 vccd1 _7409_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3055_ _6195_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3055_/X sky130_fd_sc_hd__clkbuf_16
X_5188_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5339_/B sky130_fd_sc_hd__clkbuf_2
X_4139_ _4400_/A _4265_/B vssd1 vssd1 vccd1 vccd1 _4155_/S sky130_fd_sc_hd__nor2_2
XFILLER_83_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3510_ _7082_/Q _3510_/B _5585_/B _5585_/C vssd1 vssd1 vccd1 vccd1 _3510_/X sky130_fd_sc_hd__or4_1
XFILLER_8_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4490_ _4211_/X _7309_/Q _4498_/S vssd1 vssd1 vccd1 vccd1 _4491_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__3095_ clkbuf_0__3095_/X vssd1 vssd1 vccd1 vccd1 _6370_/A sky130_fd_sc_hd__clkbuf_16
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _6462_/A _7652_/Q vssd1 vssd1 vccd1 vccd1 _6161_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5592_/D _5591_/B _7010_/A _5440_/A vssd1 vssd1 vccd1 vccd1 _5112_/A sky130_fd_sc_hd__and4_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6127_/B vssd1 vssd1 vccd1 vccd1 _6446_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5042_ _5042_/A _5046_/B vssd1 vssd1 vccd1 vccd1 _5043_/A sky130_fd_sc_hd__and2_1
XFILLER_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6993_ _6993_/A vssd1 vssd1 vccd1 vccd1 _7031_/A sky130_fd_sc_hd__clkbuf_1
X_5944_ _7396_/Q _7238_/Q _7554_/Q _7460_/Q _5921_/X _4468_/A vssd1 vssd1 vccd1 vccd1
+ _5945_/B sky130_fd_sc_hd__mux4_1
X_5875_ _5899_/S _5875_/B vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__or2_1
XFILLER_21_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7614_ _7614_/CLK _7614_/D vssd1 vssd1 vccd1 vccd1 _7614_/Q sky130_fd_sc_hd__dfxtp_1
X_4826_ _4825_/X _7128_/Q _4835_/S vssd1 vssd1 vccd1 vccd1 _4827_/A sky130_fd_sc_hd__mux2_1
X_7545_ _7545_/CLK _7545_/D vssd1 vssd1 vccd1 vccd1 _7545_/Q sky130_fd_sc_hd__dfxtp_2
X_4757_ _4757_/A vssd1 vssd1 vccd1 vccd1 _7159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4688_ _3810_/X _7213_/Q _4688_/S vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__mux2_1
X_7476_ _7476_/CLK _7476_/D vssd1 vssd1 vccd1 vccd1 _7476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3708_ _3708_/A vssd1 vssd1 vccd1 vccd1 _7630_/D sky130_fd_sc_hd__clkbuf_1
X_6427_ _6427_/A vssd1 vssd1 vccd1 vccd1 _6427_/X sky130_fd_sc_hd__buf_1
X_3639_ _4846_/A _4900_/A vssd1 vssd1 vccd1 vccd1 _3669_/S sky130_fd_sc_hd__or2_2
XFILLER_108_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6358_ _6382_/A vssd1 vssd1 vccd1 vccd1 _6358_/X sky130_fd_sc_hd__buf_1
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5309_ _6236_/C _5339_/B _5469_/C vssd1 vssd1 vccd1 vccd1 _5309_/X sky130_fd_sc_hd__a21o_1
X_5677__235 _5679__237/A vssd1 vssd1 vccd1 vccd1 _7129_/CLK sky130_fd_sc_hd__inv_2
X_6289_ _6289_/A vssd1 vssd1 vccd1 vccd1 _6289_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3107_ _6419_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3107_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6202__380 _6204__382/A vssd1 vssd1 vccd1 vccd1 _7310_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3990_ _3648_/X _7522_/Q _3994_/S vssd1 vssd1 vccd1 vccd1 _3991_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2664_ clkbuf_0__2664_/X vssd1 vssd1 vccd1 vccd1 _5578__209/A sky130_fd_sc_hd__clkbuf_16
X_4611_ _4611_/A vssd1 vssd1 vccd1 vccd1 _7256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5591_ _5592_/D _5591_/B _5591_/C vssd1 vssd1 vccd1 vccd1 _5643_/B sky130_fd_sc_hd__and3_1
X_4542_ _6236_/B _4542_/B _4606_/B vssd1 vssd1 vccd1 vccd1 _4558_/S sky130_fd_sc_hd__and3_2
X_7330_ _7674_/CLK _7330_/D vssd1 vssd1 vccd1 vccd1 _7330_/Q sky130_fd_sc_hd__dfxtp_1
X_7261_ _7261_/CLK _7261_/D vssd1 vssd1 vccd1 vccd1 _7261_/Q sky130_fd_sc_hd__dfxtp_1
X_4473_ _4473_/A _4473_/B vssd1 vssd1 vccd1 vccd1 _4474_/C sky130_fd_sc_hd__or2_1
X_7192_ _7722_/CLK _7192_/D vssd1 vssd1 vccd1 vccd1 _7192_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__3078_ clkbuf_0__3078_/X vssd1 vssd1 vccd1 vccd1 _6276__419/A sky130_fd_sc_hd__clkbuf_16
X_6143_ _6143_/A _6143_/B vssd1 vssd1 vccd1 vccd1 _6143_/Y sky130_fd_sc_hd__nor2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6074_ _7275_/Q _5748_/A _6076_/S vssd1 vssd1 vccd1 vccd1 _6075_/A sky130_fd_sc_hd__mux2_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5025_/A vssd1 vssd1 vccd1 vccd1 _5025_/X sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_17 _5995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_28 _7042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_39 _6908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6976_ _5590_/A _6976_/B vssd1 vssd1 vccd1 vccd1 _6977_/A sky130_fd_sc_hd__and2b_1
X_5927_ _5966_/A _5927_/B vssd1 vssd1 vccd1 vccd1 _5927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6655__103 _6655__103/A vssd1 vssd1 vccd1 vccd1 _7547_/CLK sky130_fd_sc_hd__inv_2
X_5858_ _7535_/Q _7676_/Q _7692_/Q _7278_/Q _5856_/X _5857_/X vssd1 vssd1 vccd1 vccd1
+ _5858_/X sky130_fd_sc_hd__mux4_2
XFILLER_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4809_ _4809_/A vssd1 vssd1 vccd1 vccd1 _7135_/D sky130_fd_sc_hd__clkbuf_1
X_5789_ _5789_/A vssd1 vssd1 vccd1 vccd1 _7203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7528_ _7528_/CLK _7528_/D vssd1 vssd1 vccd1 vccd1 _7528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7459_ _7459_/CLK _7459_/D vssd1 vssd1 vccd1 vccd1 _7459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6267__414 _6267__414/A vssd1 vssd1 vccd1 vccd1 _7354_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__3422_ clkbuf_0__3422_/X vssd1 vssd1 vccd1 vccd1 _6968__54/A sky130_fd_sc_hd__clkbuf_16
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3284_ clkbuf_0__3284_/X vssd1 vssd1 vccd1 vccd1 _6716__152/A sky130_fd_sc_hd__clkbuf_16
XFILLER_40_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6648__97 _6650__99/A vssd1 vssd1 vccd1 vccd1 _7541_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6830_ _6833_/C _6829_/C _7645_/Q vssd1 vssd1 vccd1 vccd1 _6831_/B sky130_fd_sc_hd__a21o_1
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2716_ clkbuf_0__2716_/X vssd1 vssd1 vccd1 vccd1 _5705__259/A sky130_fd_sc_hd__clkbuf_16
XFILLER_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3973_ _3652_/X _7530_/Q _3975_/S vssd1 vssd1 vccd1 vccd1 _3974_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5643_ _6234_/B _5643_/B vssd1 vssd1 vccd1 vccd1 _5647_/B sky130_fd_sc_hd__nor2_1
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5747__291 _5803__293/A vssd1 vssd1 vccd1 vccd1 _7185_/CLK sky130_fd_sc_hd__inv_2
X_7313_ _7313_/CLK _7313_/D vssd1 vssd1 vccd1 vccd1 _7313_/Q sky130_fd_sc_hd__dfxtp_1
X_4525_ _4540_/S vssd1 vssd1 vccd1 vccd1 _4534_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_116_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7244_ _7244_/CLK _7244_/D vssd1 vssd1 vccd1 vccd1 _7244_/Q sky130_fd_sc_hd__dfxtp_1
X_4456_ _5917_/A vssd1 vssd1 vccd1 vccd1 _4473_/A sky130_fd_sc_hd__clkbuf_2
X_7175_ _7175_/CLK _7175_/D vssd1 vssd1 vccd1 vccd1 _7175_/Q sky130_fd_sc_hd__dfxtp_1
X_4387_ _5337_/A _4388_/B _4386_/Y vssd1 vssd1 vccd1 vccd1 _7351_/D sky130_fd_sc_hd__o21a_1
XFILLER_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6126_ _6452_/A _6452_/B _6821_/A vssd1 vssd1 vccd1 vccd1 _6126_/Y sky130_fd_sc_hd__a21oi_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6071__347 _6071__347/A vssd1 vssd1 vccd1 vccd1 _7273_/CLK sky130_fd_sc_hd__inv_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _5008_/A _5012_/B vssd1 vssd1 vccd1 vccd1 _5009_/A sky130_fd_sc_hd__and2_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6280__422 _6281__423/A vssd1 vssd1 vccd1 vccd1 _7364_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__3267_ clkbuf_0__3267_/X vssd1 vssd1 vccd1 vccd1 _6645_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_9_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5290_ _7157_/Q _7149_/Q _5290_/S vssd1 vssd1 vccd1 vccd1 _5291_/B sky130_fd_sc_hd__mux2_1
X_4310_ _4223_/X _7372_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4311_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4241_ _4238_/X _7399_/Q _4253_/S vssd1 vssd1 vccd1 vccd1 _4242_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4172_ _4172_/A vssd1 vssd1 vccd1 vccd1 _7425_/D sky130_fd_sc_hd__clkbuf_1
X_6215__390 _6241__394/A vssd1 vssd1 vccd1 vccd1 _7320_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6813_ _6868_/A _6816_/B _6813_/C vssd1 vssd1 vccd1 vccd1 _6814_/A sky130_fd_sc_hd__and3_1
X_6744_ _6744_/A vssd1 vssd1 vccd1 vccd1 _6744_/X sky130_fd_sc_hd__buf_1
X_3956_ _3956_/A vssd1 vssd1 vccd1 vccd1 _7538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3887_ _7563_/Q _3588_/X _3891_/S vssd1 vssd1 vccd1 vccd1 _3888_/A sky130_fd_sc_hd__mux2_1
X_5626_ _5637_/A vssd1 vssd1 vccd1 vccd1 _5635_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5557_ _5444_/X _5554_/Y _5591_/C _7105_/D vssd1 vssd1 vccd1 vccd1 _5557_/X sky130_fd_sc_hd__a31o_1
XFILLER_117_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4508_ _7301_/Q _4320_/X _4516_/S vssd1 vssd1 vccd1 vccd1 _4509_/A sky130_fd_sc_hd__mux2_1
X_5488_ _5375_/X _7206_/Q input23/X _5376_/X vssd1 vssd1 vccd1 vccd1 _5488_/X sky130_fd_sc_hd__a22o_1
X_7227_ _7227_/CLK _7227_/D vssd1 vssd1 vccd1 vccd1 _7227_/Q sky130_fd_sc_hd__dfxtp_1
X_4439_ _7320_/Q _7329_/Q _4437_/Y _4438_/X vssd1 vssd1 vccd1 vccd1 _7320_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_0__3286_ _6720_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3286_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7158_ _7158_/CLK _7158_/D vssd1 vssd1 vccd1 vccd1 _7158_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _7359_/CLK _7089_/D vssd1 vssd1 vccd1 vccd1 _7089_/Q sky130_fd_sc_hd__dfxtp_2
X_6109_ _6446_/A _6127_/C _6159_/C _6109_/D vssd1 vssd1 vccd1 vccd1 _6458_/B sky130_fd_sc_hd__nor4_2
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6344__474 _6344__474/A vssd1 vssd1 vccd1 vccd1 _7416_/CLK sky130_fd_sc_hd__inv_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__3052_ clkbuf_0__3052_/X vssd1 vssd1 vccd1 vccd1 _6180__362/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6668__113 _6669__114/A vssd1 vssd1 vccd1 vccd1 _7557_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6386__508 _6387__509/A vssd1 vssd1 vccd1 vccd1 _7450_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3810_ _7670_/Q vssd1 vssd1 vccd1 vccd1 _3810_/X sky130_fd_sc_hd__buf_4
X_4790_ _7143_/Q _4569_/A _4794_/S vssd1 vssd1 vccd1 vccd1 _4791_/A sky130_fd_sc_hd__mux2_1
X_3741_ _3911_/A vssd1 vssd1 vccd1 vccd1 _3741_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6022__308 _6023__309/A vssd1 vssd1 vccd1 vccd1 _7234_/CLK sky130_fd_sc_hd__inv_2
X_3672_ _4936_/A _4542_/B vssd1 vssd1 vccd1 vccd1 _3688_/S sky130_fd_sc_hd__nand2_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6460_ _6460_/A _6509_/A vssd1 vssd1 vccd1 vccd1 _6572_/B sky130_fd_sc_hd__nor2_1
X_5411_ _5375_/X _7067_/Q _5376_/X input31/X _5410_/X vssd1 vssd1 vccd1 vccd1 _5411_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput103 _5089_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[19] sky130_fd_sc_hd__buf_2
Xoutput125 _5002_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[12] sky130_fd_sc_hd__buf_2
Xoutput114 _5054_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[3] sky130_fd_sc_hd__buf_2
X_5342_ _5236_/X _5338_/X _5339_/Y _5341_/Y vssd1 vssd1 vccd1 vccd1 _5343_/B sky130_fd_sc_hd__a31o_1
Xoutput136 _5025_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput158 _4961_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_stb_o sky130_fd_sc_hd__buf_2
Xoutput147 _4983_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[3] sky130_fd_sc_hd__buf_2
Xoutput169 _5473_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[17] sky130_fd_sc_hd__buf_2
X_7012_ _6923_/A _6476_/A _7024_/S vssd1 vssd1 vccd1 vccd1 _7013_/B sky130_fd_sc_hd__mux2_1
X_5273_ _5264_/X _5266_/Y _5269_/X _5272_/Y vssd1 vssd1 vccd1 vccd1 _5273_/X sky130_fd_sc_hd__a31o_1
XFILLER_101_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4224_ _4223_/X _7404_/Q _4227_/S vssd1 vssd1 vccd1 vccd1 _4225_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4155_ _7432_/Q _3603_/X _4155_/S vssd1 vssd1 vccd1 vccd1 _4156_/A sky130_fd_sc_hd__mux2_1
X_6287__428 _6287__428/A vssd1 vssd1 vccd1 vccd1 _7370_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4086_ _7459_/Q _3810_/X _4086_/S vssd1 vssd1 vccd1 vccd1 _4087_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4988_ _6921_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__and2_1
X_3939_ _3656_/X _7545_/Q _3939_/S vssd1 vssd1 vccd1 vccd1 _3940_/A sky130_fd_sc_hd__mux2_1
X_6658_ _6664_/A vssd1 vssd1 vccd1 vccd1 _6658_/X sky130_fd_sc_hd__buf_1
X_5609_ _7088_/Q _5066_/A _5613_/S vssd1 vssd1 vccd1 vccd1 _5610_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6589_ _7509_/Q _6589_/B _6594_/C vssd1 vssd1 vccd1 vccd1 _6589_/X sky130_fd_sc_hd__and3_1
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3269_ _6633_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3269_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3104_ clkbuf_0__3104_/X vssd1 vssd1 vccd1 vccd1 _6406__524/A sky130_fd_sc_hd__clkbuf_16
Xinput16 caravel_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_2
Xinput27 caravel_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_2
X_6392__512 _6392__512/A vssd1 vssd1 vccd1 vccd1 _7454_/CLK sky130_fd_sc_hd__inv_2
Xinput38 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 _5068_/A sky130_fd_sc_hd__buf_4
Xinput49 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _5060_/A sky130_fd_sc_hd__buf_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5960_ _5956_/X _5959_/X _5999_/S vssd1 vssd1 vccd1 vccd1 _5960_/X sky130_fd_sc_hd__mux2_2
XFILLER_65_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5891_ _7410_/Q _7378_/Q _7709_/Q _7632_/Q _5857_/X _4484_/X vssd1 vssd1 vccd1 vccd1
+ _5891_/X sky130_fd_sc_hd__mux4_1
X_4911_ _4911_/A vssd1 vssd1 vccd1 vccd1 _7056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5670__230 _5674__234/A vssd1 vssd1 vccd1 vccd1 _7124_/CLK sky130_fd_sc_hd__inv_2
X_7630_ _7630_/CLK _7630_/D vssd1 vssd1 vccd1 vccd1 _7630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4842_ _4842_/A vssd1 vssd1 vccd1 vccd1 _7123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7561_ _7561_/CLK _7561_/D vssd1 vssd1 vccd1 vccd1 _7561_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4773_ _4773_/A vssd1 vssd1 vccd1 vccd1 _7151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3724_ _3538_/X _7624_/Q _3728_/S vssd1 vssd1 vccd1 vccd1 _3725_/A sky130_fd_sc_hd__mux2_1
X_7492_ _7492_/CLK _7492_/D vssd1 vssd1 vccd1 vccd1 _7492_/Q sky130_fd_sc_hd__dfxtp_1
X_6512_ _6525_/A vssd1 vssd1 vccd1 vccd1 _6534_/A sky130_fd_sc_hd__clkbuf_2
X_3655_ _7324_/Q vssd1 vssd1 vccd1 vccd1 _4575_/A sky130_fd_sc_hd__clkbuf_4
X_3586_ _7705_/Q _3585_/X _3595_/S vssd1 vssd1 vccd1 vccd1 _3587_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5325_ _7290_/Q _7703_/Q _5325_/S vssd1 vssd1 vccd1 vccd1 _5325_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5256_ _7528_/Q _7108_/Q _7560_/Q _7124_/Q _5132_/X _5135_/X vssd1 vssd1 vccd1 vccd1
+ _5257_/B sky130_fd_sc_hd__mux4_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4207_ _4115_/X _7409_/Q _4209_/S vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3054_ _6189_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3054_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5187_ _5187_/A _5380_/C _5187_/C vssd1 vssd1 vccd1 vccd1 _5188_/A sky130_fd_sc_hd__nor3_1
XFILLER_110_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4138_ _4138_/A vssd1 vssd1 vccd1 vccd1 _7440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4069_ _4069_/A vssd1 vssd1 vccd1 vccd1 _7467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6194__374 _6194__374/A vssd1 vssd1 vccd1 vccd1 _7304_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5734__282 _5735__283/A vssd1 vssd1 vccd1 vccd1 _7176_/CLK sky130_fd_sc_hd__inv_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__3094_ clkbuf_0__3094_/X vssd1 vssd1 vccd1 vccd1 _6355__483/A sky130_fd_sc_hd__clkbuf_16
XFILLER_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5741__286 _5743__288/A vssd1 vssd1 vccd1 vccd1 _7180_/CLK sky130_fd_sc_hd__inv_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5185_/B vssd1 vssd1 vccd1 vccd1 _5440_/A sky130_fd_sc_hd__clkbuf_2
X_6090_ _7731_/Q _7730_/Q _7729_/Q _7728_/Q vssd1 vssd1 vccd1 vccd1 _6127_/B sky130_fd_sc_hd__or4_1
X_5041_ _5041_/A vssd1 vssd1 vccd1 vccd1 _5041_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_6992_ _6992_/A vssd1 vssd1 vccd1 vccd1 _7719_/D sky130_fd_sc_hd__clkbuf_1
X_5943_ _6005_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6399__518 _6399__518/A vssd1 vssd1 vccd1 vccd1 _7460_/CLK sky130_fd_sc_hd__inv_2
X_5874_ _7409_/Q _7377_/Q _7708_/Q _7631_/Q _5921_/A _5818_/X vssd1 vssd1 vccd1 vccd1
+ _5875_/B sky130_fd_sc_hd__mux4_1
XFILLER_80_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7613_ _7613_/CLK _7613_/D vssd1 vssd1 vccd1 vccd1 _7613_/Q sky130_fd_sc_hd__dfxtp_2
X_4825_ _7327_/Q vssd1 vssd1 vccd1 vccd1 _4825_/X sky130_fd_sc_hd__buf_2
X_7544_ _7544_/CLK _7544_/D vssd1 vssd1 vccd1 vccd1 _7544_/Q sky130_fd_sc_hd__dfxtp_1
X_4756_ _4569_/X _7159_/Q _4760_/S vssd1 vssd1 vccd1 vccd1 _4757_/A sky130_fd_sc_hd__mux2_1
X_7475_ _7475_/CLK _7475_/D vssd1 vssd1 vccd1 vccd1 _7475_/Q sky130_fd_sc_hd__dfxtp_1
X_4687_ _4687_/A vssd1 vssd1 vccd1 vccd1 _7214_/D sky130_fd_sc_hd__clkbuf_1
X_3707_ _3546_/X _7630_/Q _3707_/S vssd1 vssd1 vccd1 vccd1 _3708_/A sky130_fd_sc_hd__mux2_1
X_3638_ _4363_/A _3927_/C _3927_/A vssd1 vssd1 vccd1 vccd1 _4900_/A sky130_fd_sc_hd__or3b_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6357_ _6357_/A vssd1 vssd1 vccd1 vccd1 _6357_/X sky130_fd_sc_hd__buf_1
X_3569_ _3756_/A _4376_/B _3560_/Y _3568_/X vssd1 vssd1 vccd1 vccd1 _3573_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_102_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5308_ _5308_/A _5308_/B _5308_/C vssd1 vssd1 vccd1 vccd1 _5308_/Y sky130_fd_sc_hd__nor3_2
Xclkbuf_0__3106_ _6413_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3106_/X sky130_fd_sc_hd__clkbuf_16
X_6035__318 _6035__318/A vssd1 vssd1 vccd1 vccd1 _7244_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5239_ _5239_/A _5239_/B vssd1 vssd1 vccd1 vccd1 _5240_/A sky130_fd_sc_hd__or2_1
XFILLER_29_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4610_ _7256_/Q _3905_/A _4616_/S vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5590_ _5590_/A _5590_/B vssd1 vssd1 vccd1 vccd1 _7080_/D sky130_fd_sc_hd__nor2_1
X_4541_ _4541_/A vssd1 vssd1 vccd1 vccd1 _7286_/D sky130_fd_sc_hd__clkbuf_1
X_7260_ _7260_/CLK _7260_/D vssd1 vssd1 vccd1 vccd1 _7260_/Q sky130_fd_sc_hd__dfxtp_1
X_4472_ _5832_/A _4474_/B _4471_/Y _4438_/X vssd1 vssd1 vccd1 vccd1 _7314_/D sky130_fd_sc_hd__o211a_1
XFILLER_7_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7191_ _7732_/CLK _7191_/D vssd1 vssd1 vccd1 vccd1 _7191_/Q sky130_fd_sc_hd__dfxtp_1
X_6142_ _7730_/Q _7641_/Q vssd1 vssd1 vccd1 vccd1 _6143_/B sky130_fd_sc_hd__xnor2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3077_ clkbuf_0__3077_/X vssd1 vssd1 vccd1 vccd1 _6267__414/A sky130_fd_sc_hd__clkbuf_16
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6073_ _6073_/A vssd1 vssd1 vccd1 vccd1 _7274_/D sky130_fd_sc_hd__clkbuf_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5024_/A _5024_/B vssd1 vssd1 vccd1 vccd1 _5025_/A sky130_fd_sc_hd__and2_1
XFILLER_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_18 _6005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_29 _7043_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6975_ _5012_/A _7715_/Q _6978_/S vssd1 vssd1 vccd1 vccd1 _6976_/B sky130_fd_sc_hd__mux2_1
X_5926_ _7625_/Q _7617_/Q _7601_/Q _7593_/Q _5870_/X _5925_/X vssd1 vssd1 vccd1 vccd1
+ _5927_/B sky130_fd_sc_hd__mux4_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5857_ _5857_/A vssd1 vssd1 vccd1 vccd1 _5857_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4808_ _4569_/X _7135_/Q _4812_/S vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__mux2_1
X_5788_ _7203_/Q _5031_/A _5794_/S vssd1 vssd1 vccd1 vccd1 _5789_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7527_ _7527_/CLK _7527_/D vssd1 vssd1 vccd1 vccd1 _7527_/Q sky130_fd_sc_hd__dfxtp_1
X_5683__240 _5686__243/A vssd1 vssd1 vccd1 vccd1 _7134_/CLK sky130_fd_sc_hd__inv_2
X_4739_ _4739_/A vssd1 vssd1 vccd1 vccd1 _7167_/D sky130_fd_sc_hd__clkbuf_1
X_7458_ _7458_/CLK _7458_/D vssd1 vssd1 vccd1 vccd1 _7458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7389_ _7389_/CLK _7389_/D vssd1 vssd1 vccd1 vccd1 _7389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6662__108 _6662__108/A vssd1 vssd1 vccd1 vccd1 _7552_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3421_ clkbuf_0__3421_/X vssd1 vssd1 vccd1 vccd1 _6961__48/A sky130_fd_sc_hd__clkbuf_16
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6424__57 _6424__57/A vssd1 vssd1 vccd1 vccd1 _7479_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3283_ clkbuf_0__3283_/X vssd1 vssd1 vccd1 vccd1 _6712__149/A sky130_fd_sc_hd__clkbuf_16
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__2715_ clkbuf_0__2715_/X vssd1 vssd1 vccd1 vccd1 _5698__253/A sky130_fd_sc_hd__clkbuf_16
X_3972_ _3972_/A vssd1 vssd1 vccd1 vccd1 _7531_/D sky130_fd_sc_hd__clkbuf_1
X_5642_ _5642_/A _6234_/B vssd1 vssd1 vccd1 vccd1 _5642_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5573_ _5573_/A vssd1 vssd1 vccd1 vccd1 _5573_/X sky130_fd_sc_hd__buf_1
XFILLER_116_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4524_ _4882_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4540_/S sky130_fd_sc_hd__or2_2
X_7312_ _7312_/CLK _7312_/D vssd1 vssd1 vccd1 vccd1 _7312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7243_ _7243_/CLK _7243_/D vssd1 vssd1 vccd1 vccd1 _7243_/Q sky130_fd_sc_hd__dfxtp_1
X_4455_ _5929_/A vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7174_ _7174_/CLK _7174_/D vssd1 vssd1 vccd1 vccd1 _7174_/Q sky130_fd_sc_hd__dfxtp_1
X_4386_ _5337_/A _4388_/B _6274_/A vssd1 vssd1 vccd1 vccd1 _4386_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6125_ _7643_/Q vssd1 vssd1 vccd1 vccd1 _6821_/A sky130_fd_sc_hd__clkbuf_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6056_/A vssd1 vssd1 vccd1 vccd1 _6056_/X sky130_fd_sc_hd__buf_1
XFILLER_65_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5007_ _5007_/A vssd1 vssd1 vccd1 vccd1 _5007_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5909_ _7585_/Q _7577_/Q _7569_/Q _7483_/Q _5907_/X _5908_/X vssd1 vssd1 vccd1 vccd1
+ _5909_/X sky130_fd_sc_hd__mux4_2
X_6889_ _6889_/A _6889_/B vssd1 vssd1 vccd1 vccd1 _6903_/B sky130_fd_sc_hd__or2_1
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6087__355 _6173__357/A vssd1 vssd1 vccd1 vccd1 _7284_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3266_ clkbuf_0__3266_/X vssd1 vssd1 vccd1 vccd1 _6621__76/A sky130_fd_sc_hd__clkbuf_16
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4240_ _4262_/S vssd1 vssd1 vccd1 vccd1 _4253_/S sky130_fd_sc_hd__buf_2
XFILLER_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4171_ _4115_/X _7425_/Q _4173_/S vssd1 vssd1 vccd1 vccd1 _4172_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6812_ _7641_/Q _6819_/D vssd1 vssd1 vccd1 vccd1 _6813_/C sky130_fd_sc_hd__or2_1
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3955_ _3911_/X _7538_/Q _3957_/S vssd1 vssd1 vccd1 vccd1 _3956_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2629_ clkbuf_0__2629_/X vssd1 vssd1 vccd1 vccd1 _5573_/A sky130_fd_sc_hd__clkbuf_16
X_3886_ _3886_/A vssd1 vssd1 vccd1 vccd1 _7564_/D sky130_fd_sc_hd__clkbuf_1
X_5625_ _5625_/A vssd1 vssd1 vccd1 vccd1 _7095_/D sky130_fd_sc_hd__clkbuf_1
X_5556_ _7070_/Q _7069_/Q _5554_/Y vssd1 vssd1 vccd1 vccd1 _7105_/D sky130_fd_sc_hd__o21a_1
X_5487_ _5481_/X _7205_/Q input22/X _5482_/X vssd1 vssd1 vccd1 vccd1 _5487_/X sky130_fd_sc_hd__a22o_2
X_4507_ _4522_/S vssd1 vssd1 vccd1 vccd1 _4516_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7226_ _7226_/CLK _7226_/D vssd1 vssd1 vccd1 vccd1 _7226_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3285_ _6719_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3285_/X sky130_fd_sc_hd__clkbuf_16
X_4438_ _6236_/B vssd1 vssd1 vccd1 vccd1 _4438_/X sky130_fd_sc_hd__buf_2
XFILLER_104_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7157_ _7157_/CLK _7157_/D vssd1 vssd1 vccd1 vccd1 _7157_/Q sky130_fd_sc_hd__dfxtp_1
X_4369_ _7349_/Q vssd1 vssd1 vccd1 vccd1 _5262_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7088_/CLK _7088_/D vssd1 vssd1 vccd1 vccd1 _7088_/Q sky130_fd_sc_hd__dfxtp_1
X_6108_ _7719_/Q _7718_/Q vssd1 vssd1 vccd1 vccd1 _6109_/D sky130_fd_sc_hd__or2_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3051_ clkbuf_0__3051_/X vssd1 vssd1 vccd1 vccd1 _6201_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6238__391 _6241__394/A vssd1 vssd1 vccd1 vccd1 _7331_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6936__28 _6937__29/A vssd1 vssd1 vccd1 vccd1 _7684_/CLK sky130_fd_sc_hd__inv_2
X_3740_ _3740_/A vssd1 vssd1 vccd1 vccd1 _7619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3671_ _3671_/A _4436_/A _3711_/C vssd1 vssd1 vccd1 vccd1 _4936_/A sky130_fd_sc_hd__and3_4
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5410_ _5494_/S _5436_/B _5410_/C vssd1 vssd1 vccd1 vccd1 _5410_/X sky130_fd_sc_hd__and3_1
Xoutput115 _5056_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[4] sky130_fd_sc_hd__buf_2
Xoutput104 _5050_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[1] sky130_fd_sc_hd__buf_2
X_5341_ _6784_/A _5236_/X _5112_/X vssd1 vssd1 vccd1 vccd1 _5341_/Y sky130_fd_sc_hd__o21ai_1
Xoutput137 _5028_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput126 _5005_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput159 _4963_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_we_o sky130_fd_sc_hd__buf_2
Xoutput148 _4985_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_99_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7011_ _7033_/S vssd1 vssd1 vccd1 vccd1 _7024_/S sky130_fd_sc_hd__clkbuf_2
X_5272_ _5349_/S _5271_/X _5178_/A vssd1 vssd1 vccd1 vccd1 _5272_/Y sky130_fd_sc_hd__o21ai_1
X_4223_ _4572_/A vssd1 vssd1 vccd1 vccd1 _4223_/X sky130_fd_sc_hd__clkbuf_4
X_4154_ _4154_/A vssd1 vssd1 vccd1 vccd1 _7433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4085_ _4085_/A vssd1 vssd1 vccd1 vccd1 _7460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4987_ _4987_/A vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__clkbuf_1
X_6726_ _6732_/A vssd1 vssd1 vccd1 vccd1 _6726_/X sky130_fd_sc_hd__buf_1
XFILLER_51_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3938_ _3938_/A vssd1 vssd1 vccd1 vccd1 _7546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3869_ _3869_/A vssd1 vssd1 vccd1 vccd1 _7571_/D sky130_fd_sc_hd__clkbuf_1
X_6657_ _6688_/A vssd1 vssd1 vccd1 vccd1 _6657_/X sky130_fd_sc_hd__buf_1
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5608_ _5608_/A vssd1 vssd1 vccd1 vccd1 _7087_/D sky130_fd_sc_hd__clkbuf_1
X_6588_ _6592_/B _6588_/B _6593_/C vssd1 vssd1 vccd1 vccd1 _6588_/X sky130_fd_sc_hd__and3b_1
X_5539_ _5539_/A vssd1 vssd1 vccd1 vccd1 _7061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3268_ _6626_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3268_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7209_ _7510_/CLK _7209_/D vssd1 vssd1 vccd1 vccd1 _7209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3103_ clkbuf_0__3103_/X vssd1 vssd1 vccd1 vccd1 _6400__519/A sky130_fd_sc_hd__clkbuf_16
XFILLER_23_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput17 caravel_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_2
Xinput28 caravel_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_4
X_6941__31 _6941__31/A vssd1 vssd1 vccd1 vccd1 _7687_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput39 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__buf_4
XFILLER_2_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5890_ _5966_/A _5890_/B vssd1 vssd1 vccd1 vccd1 _5890_/Y sky130_fd_sc_hd__nor2_1
X_4910_ _4834_/X _7056_/Q _4910_/S vssd1 vssd1 vccd1 vccd1 _4911_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4841_ _4840_/X _7123_/Q _4844_/S vssd1 vssd1 vccd1 vccd1 _4842_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7560_ _7560_/CLK _7560_/D vssd1 vssd1 vccd1 vccd1 _7560_/Q sky130_fd_sc_hd__dfxtp_2
X_4772_ _7151_/Q _4328_/X _4774_/S vssd1 vssd1 vccd1 vccd1 _4773_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3723_ _3723_/A vssd1 vssd1 vccd1 vccd1 _7625_/D sky130_fd_sc_hd__clkbuf_1
X_7491_ _7491_/CLK _7491_/D vssd1 vssd1 vccd1 vccd1 _7491_/Q sky130_fd_sc_hd__dfxtp_1
X_6511_ _6504_/X _6460_/A _6509_/X _6510_/X vssd1 vssd1 vccd1 vccd1 _6525_/A sky130_fd_sc_hd__o31a_1
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3654_ _3654_/A vssd1 vssd1 vccd1 vccd1 _7687_/D sky130_fd_sc_hd__clkbuf_1
X_6293__433 _6294__434/A vssd1 vssd1 vccd1 vccd1 _7375_/CLK sky130_fd_sc_hd__inv_2
X_3585_ _7327_/Q vssd1 vssd1 vccd1 vccd1 _3585_/X sky130_fd_sc_hd__buf_4
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5324_ _5331_/A _5324_/B vssd1 vssd1 vccd1 vccd1 _5324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5255_ _5205_/X _5248_/X _5250_/Y _5254_/Y vssd1 vssd1 vccd1 vccd1 _5255_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_114_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4206_ _4206_/A vssd1 vssd1 vccd1 vccd1 _7410_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3053_ _6183_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3053_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5186_ _5585_/B _5440_/A _5232_/A _5185_/Y _7081_/Q vssd1 vssd1 vccd1 vccd1 _5187_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _4118_/X _7440_/Q _4137_/S vssd1 vssd1 vccd1 vccd1 _4138_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4068_ _3914_/X _7467_/Q _4068_/S vssd1 vssd1 vccd1 vccd1 _4069_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7689_ _7689_/CLK _7689_/D vssd1 vssd1 vccd1 vccd1 _7689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3093_ clkbuf_0__3093_/X vssd1 vssd1 vccd1 vccd1 _6347__476/A sky130_fd_sc_hd__clkbuf_16
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/A _5046_/B vssd1 vssd1 vccd1 vccd1 _5041_/A sky130_fd_sc_hd__and2_1
XFILLER_111_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6991_ _6981_/X _6991_/B vssd1 vssd1 vccd1 vccd1 _6992_/A sky130_fd_sc_hd__and2b_1
XFILLER_26_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5942_ _7452_/Q _7444_/Q _7428_/Q _7420_/Q _5856_/X _5857_/X vssd1 vssd1 vccd1 vccd1
+ _5943_/B sky130_fd_sc_hd__mux4_1
XFILLER_65_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5873_ _7623_/Q _7615_/Q _7599_/Q _7591_/Q _5851_/X _5852_/X vssd1 vssd1 vccd1 vccd1
+ _5873_/X sky130_fd_sc_hd__mux4_2
X_7612_ _7612_/CLK _7612_/D vssd1 vssd1 vccd1 vccd1 _7612_/Q sky130_fd_sc_hd__dfxtp_2
X_4824_ _4824_/A vssd1 vssd1 vccd1 vccd1 _7129_/D sky130_fd_sc_hd__clkbuf_1
X_7543_ _7543_/CLK _7543_/D vssd1 vssd1 vccd1 vccd1 _7543_/Q sky130_fd_sc_hd__dfxtp_2
X_4755_ _4755_/A vssd1 vssd1 vccd1 vccd1 _7160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3706_ _3706_/A vssd1 vssd1 vccd1 vccd1 _7631_/D sky130_fd_sc_hd__clkbuf_1
X_4686_ _3807_/X _7214_/Q _4688_/S vssd1 vssd1 vccd1 vccd1 _4687_/A sky130_fd_sc_hd__mux2_1
X_7474_ _7474_/CLK _7474_/D vssd1 vssd1 vccd1 vccd1 _7474_/Q sky130_fd_sc_hd__dfxtp_1
X_3637_ _4363_/B _6222_/A vssd1 vssd1 vccd1 vccd1 _3927_/C sky130_fd_sc_hd__nand2_1
XFILLER_115_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3568_ _7347_/Q _3570_/C vssd1 vssd1 vccd1 vccd1 _3568_/X sky130_fd_sc_hd__and2b_1
XFILLER_103_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5307_ _5131_/X _5301_/X _5306_/X _5161_/X vssd1 vssd1 vccd1 vccd1 _5308_/C sky130_fd_sc_hd__a211oi_1
Xclkbuf_0__3105_ _6407_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3105_/X sky130_fd_sc_hd__clkbuf_16
X_3499_ _7103_/Q vssd1 vssd1 vccd1 vccd1 _6910_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5238_ _5238_/A _5238_/B vssd1 vssd1 vccd1 vccd1 _5239_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5169_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5173_/A sky130_fd_sc_hd__buf_2
XFILLER_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _4235_/X _7286_/Q _4540_/S vssd1 vssd1 vccd1 vccd1 _4541_/A sky130_fd_sc_hd__mux2_1
X_4471_ _5832_/A _4474_/B vssd1 vssd1 vccd1 vccd1 _4471_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7190_ _7190_/CLK _7190_/D vssd1 vssd1 vccd1 vccd1 _7190_/Q sky130_fd_sc_hd__dfxtp_1
X_6141_ _6487_/A _7640_/Q vssd1 vssd1 vccd1 vccd1 _6143_/A sky130_fd_sc_hd__and2b_1
Xclkbuf_1_0__f__3076_ clkbuf_0__3076_/X vssd1 vssd1 vccd1 vccd1 _6277_/A sky130_fd_sc_hd__clkbuf_16
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6072_ _7010_/A _5536_/A _6076_/S vssd1 vssd1 vccd1 vccd1 _6073_/A sky130_fd_sc_hd__mux2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5023_/A vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_19 _7304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6974_ _7276_/Q _7010_/B vssd1 vssd1 vccd1 vccd1 _6978_/S sky130_fd_sc_hd__nand2_1
XFILLER_110_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5925_ _5925_/A vssd1 vssd1 vccd1 vccd1 _5925_/X sky130_fd_sc_hd__clkbuf_2
X_5856_ _5856_/A vssd1 vssd1 vccd1 vccd1 _5856_/X sky130_fd_sc_hd__buf_4
X_4807_ _4807_/A vssd1 vssd1 vccd1 vccd1 _7136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6041__323 _6041__323/A vssd1 vssd1 vccd1 vccd1 _7249_/CLK sky130_fd_sc_hd__inv_2
X_5787_ _5787_/A vssd1 vssd1 vccd1 vccd1 _7202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7526_ _7526_/CLK _7526_/D vssd1 vssd1 vccd1 vccd1 _7526_/Q sky130_fd_sc_hd__dfxtp_1
X_4738_ _7167_/Q _4328_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4739_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4669_ _4669_/A vssd1 vssd1 vccd1 vccd1 _7230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7457_ _7457_/CLK _7457_/D vssd1 vssd1 vccd1 vccd1 _7457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7388_ _7388_/CLK _7388_/D vssd1 vssd1 vccd1 vccd1 _7388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6339_ _6351_/A vssd1 vssd1 vccd1 vccd1 _6339_/X sky130_fd_sc_hd__buf_1
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3420_ clkbuf_0__3420_/X vssd1 vssd1 vccd1 vccd1 _6955__43/A sky130_fd_sc_hd__clkbuf_16
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__3282_ clkbuf_0__3282_/X vssd1 vssd1 vccd1 vccd1 _6706__144/A sky130_fd_sc_hd__clkbuf_16
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3971_ _3648_/X _7531_/Q _3975_/S vssd1 vssd1 vccd1 vccd1 _3972_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2714_ clkbuf_0__2714_/X vssd1 vssd1 vccd1 vccd1 _5693__249/A sky130_fd_sc_hd__clkbuf_16
XFILLER_16_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5641_ _5641_/A vssd1 vssd1 vccd1 vccd1 _7102_/D sky130_fd_sc_hd__clkbuf_1
X_7311_ _7311_/CLK _7311_/D vssd1 vssd1 vccd1 vccd1 _7311_/Q sky130_fd_sc_hd__dfxtp_2
X_4523_ _4523_/A vssd1 vssd1 vccd1 vccd1 _7294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7242_ _7242_/CLK _7242_/D vssd1 vssd1 vccd1 vccd1 _7242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4454_ _7314_/Q vssd1 vssd1 vccd1 vccd1 _5832_/A sky130_fd_sc_hd__inv_2
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7173_ _7173_/CLK _7173_/D vssd1 vssd1 vccd1 vccd1 _7173_/Q sky130_fd_sc_hd__dfxtp_1
X_4385_ _4385_/A vssd1 vssd1 vccd1 vccd1 _6274_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6124_ _5235_/X _6119_/B _7729_/Q _6784_/A vssd1 vssd1 vccd1 vccd1 _6452_/B sky130_fd_sc_hd__o31ai_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3059_ clkbuf_0__3059_/X vssd1 vssd1 vccd1 vccd1 _6241__394/A sky130_fd_sc_hd__clkbuf_16
XFILLER_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6055_ _6055_/A vssd1 vssd1 vccd1 vccd1 _6055_/X sky130_fd_sc_hd__buf_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5006_/A _5012_/B vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__and2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _6963_/A vssd1 vssd1 vccd1 vccd1 _6957_/X sky130_fd_sc_hd__buf_1
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5908_ _5908_/A vssd1 vssd1 vccd1 vccd1 _5908_/X sky130_fd_sc_hd__clkbuf_2
X_6888_ _6794_/A _6781_/X _6886_/X _6887_/X vssd1 vssd1 vccd1 vccd1 _7658_/D sky130_fd_sc_hd__o211a_1
X_5839_ _5855_/A vssd1 vssd1 vccd1 vccd1 _5910_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7509_ _7510_/CLK _7509_/D vssd1 vssd1 vccd1 vccd1 _7509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6048__329 _6048__329/A vssd1 vssd1 vccd1 vccd1 _7255_/CLK sky130_fd_sc_hd__inv_2
X_6948__37 _6948__37/A vssd1 vssd1 vccd1 vccd1 _7693_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _4170_/A vssd1 vssd1 vccd1 vccd1 _7426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6811_ _7641_/Q _6819_/D vssd1 vssd1 vccd1 vccd1 _6816_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3954_ _3954_/A vssd1 vssd1 vccd1 vccd1 _7539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3885_ _7564_/Q _3585_/X _3891_/S vssd1 vssd1 vccd1 vccd1 _3886_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__2628_ clkbuf_0__2628_/X vssd1 vssd1 vccd1 vccd1 _5504__184/A sky130_fd_sc_hd__clkbuf_16
XFILLER_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5624_ _7095_/Q _7194_/Q _5624_/S vssd1 vssd1 vccd1 vccd1 _5625_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3422_ _6963_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3422_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5555_ _5555_/A _5555_/B vssd1 vssd1 vccd1 vccd1 _5591_/C sky130_fd_sc_hd__and2_2
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5486_ _5481_/X _7204_/Q input21/X _5482_/X vssd1 vssd1 vccd1 vccd1 _5486_/X sky130_fd_sc_hd__a22o_2
X_4506_ _4562_/A _4506_/B vssd1 vssd1 vccd1 vccd1 _4522_/S sky130_fd_sc_hd__nor2_2
Xclkbuf_0__3284_ _6713_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3284_/X sky130_fd_sc_hd__clkbuf_16
X_7225_ _7516_/CLK _7225_/D vssd1 vssd1 vccd1 vccd1 _7225_/Q sky130_fd_sc_hd__dfxtp_1
X_4437_ _4443_/B vssd1 vssd1 vccd1 vccd1 _4437_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7156_ _7156_/CLK _7156_/D vssd1 vssd1 vccd1 vccd1 _7156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _6107_/A _6792_/B vssd1 vssd1 vccd1 vccd1 _6778_/B sky130_fd_sc_hd__xor2_1
X_4368_ _4368_/A vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4299_ _4261_/X _7376_/Q _4299_/S vssd1 vssd1 vccd1 vccd1 _4300_/A sky130_fd_sc_hd__mux2_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _7359_/CLK _7087_/D vssd1 vssd1 vccd1 vccd1 _7087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5696__251 _5698__253/A vssd1 vssd1 vccd1 vccd1 _7145_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7190_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6675__119 _6675__119/A vssd1 vssd1 vccd1 vccd1 _7563_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3670_ _3670_/A vssd1 vssd1 vccd1 vccd1 _7683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput105 _5091_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput116 _5058_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[5] sky130_fd_sc_hd__buf_2
XFILLER_114_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5340_ _7728_/Q vssd1 vssd1 vccd1 vccd1 _6784_/A sky130_fd_sc_hd__clkbuf_4
Xoutput138 _5030_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput127 _5007_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput149 _4987_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5271_ _7172_/Q _7304_/Q _7490_/Q _7180_/Q _5207_/A _5290_/S vssd1 vssd1 vccd1 vccd1
+ _5271_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4222_ _4222_/A vssd1 vssd1 vccd1 vccd1 _7405_/D sky130_fd_sc_hd__clkbuf_1
X_7010_ _7010_/A _7010_/B vssd1 vssd1 vccd1 vccd1 _7033_/S sky130_fd_sc_hd__nand2_2
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4153_ _7433_/Q _3600_/X _4155_/S vssd1 vssd1 vccd1 vccd1 _4154_/A sky130_fd_sc_hd__mux2_1
X_4084_ _7460_/Q _3807_/X _4086_/S vssd1 vssd1 vccd1 vccd1 _4085_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4986_ _6919_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4987_/A sky130_fd_sc_hd__and2_1
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3937_ _3652_/X _7546_/Q _3939_/S vssd1 vssd1 vccd1 vccd1 _3938_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3868_ _3738_/X _7571_/Q _3872_/S vssd1 vssd1 vccd1 vccd1 _3869_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3799_ _7597_/Q _3794_/X _3811_/S vssd1 vssd1 vccd1 vccd1 _3800_/A sky130_fd_sc_hd__mux2_1
X_5607_ _7087_/Q _5064_/A _5613_/S vssd1 vssd1 vccd1 vccd1 _5608_/A sky130_fd_sc_hd__mux2_1
X_6587_ _7509_/Q _6587_/B vssd1 vssd1 vccd1 vccd1 _6588_/B sky130_fd_sc_hd__or2_1
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5538_ _6908_/A _7061_/Q _5546_/S vssd1 vssd1 vccd1 vccd1 _5539_/A sky130_fd_sc_hd__mux2_1
X_5469_ _5469_/A _7276_/Q _5469_/C vssd1 vssd1 vccd1 vccd1 _5469_/X sky130_fd_sc_hd__and3_1
X_7208_ _7510_/CLK _7208_/D vssd1 vssd1 vccd1 vccd1 _7208_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3267_ _6625_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3267_/X sky130_fd_sc_hd__clkbuf_16
X_7139_ _7139_/CLK _7139_/D vssd1 vssd1 vccd1 vccd1 _7139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3102_ clkbuf_0__3102_/X vssd1 vssd1 vccd1 vccd1 _6392__512/A sky130_fd_sc_hd__clkbuf_16
Xinput18 caravel_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_2
Xinput29 caravel_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2962_ clkbuf_0__2962_/X vssd1 vssd1 vccd1 vccd1 _6071__347/A sky130_fd_sc_hd__clkbuf_16
XFILLER_38_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4840_ _7322_/Q vssd1 vssd1 vccd1 vccd1 _4840_/X sky130_fd_sc_hd__buf_2
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _4771_/A vssd1 vssd1 vccd1 vccd1 _7152_/D sky130_fd_sc_hd__clkbuf_1
X_6510_ _7497_/Q _7496_/Q vssd1 vssd1 vccd1 vccd1 _6510_/X sky130_fd_sc_hd__or2_1
X_3722_ _3534_/X _7625_/Q _3722_/S vssd1 vssd1 vccd1 vccd1 _3723_/A sky130_fd_sc_hd__mux2_1
X_7490_ _7490_/CLK _7490_/D vssd1 vssd1 vccd1 vccd1 _7490_/Q sky130_fd_sc_hd__dfxtp_1
X_3653_ _3652_/X _7687_/Q _3657_/S vssd1 vssd1 vccd1 vccd1 _3654_/A sky130_fd_sc_hd__mux2_1
X_3584_ _3584_/A vssd1 vssd1 vccd1 vccd1 _7706_/D sky130_fd_sc_hd__clkbuf_1
X_5323_ _7076_/Q _7364_/Q _5330_/S vssd1 vssd1 vccd1 vccd1 _5324_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5254_ _5356_/A _5253_/X _5178_/X vssd1 vssd1 vccd1 vccd1 _5254_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_102_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4205_ _4112_/X _7410_/Q _4209_/S vssd1 vssd1 vccd1 vccd1 _4206_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3052_ _6177_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3052_/X sky130_fd_sc_hd__clkbuf_16
X_5185_ _7082_/Q _5185_/B vssd1 vssd1 vccd1 vccd1 _5185_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4136_ _4136_/A vssd1 vssd1 vccd1 vccd1 _7441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ _4067_/A vssd1 vssd1 vccd1 vccd1 _7468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6620__75 _6621__76/A vssd1 vssd1 vccd1 vccd1 _7518_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4969_ _5106_/B vssd1 vssd1 vccd1 vccd1 _4979_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7688_ _7688_/CLK _7688_/D vssd1 vssd1 vccd1 vccd1 _7688_/Q sky130_fd_sc_hd__dfxtp_1
X_6639_ _6645_/A vssd1 vssd1 vccd1 vccd1 _6639_/X sky130_fd_sc_hd__buf_1
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6745__175 _6749__179/A vssd1 vssd1 vccd1 vccd1 _7619_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__3092_ clkbuf_0__3092_/X vssd1 vssd1 vccd1 vccd1 _6344__474/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6990_ _5004_/A _6462_/A _7000_/S vssd1 vssd1 vccd1 vccd1 _6991_/B sky130_fd_sc_hd__mux2_1
X_5941_ _5937_/X _5940_/X _5999_/S vssd1 vssd1 vccd1 vccd1 _5941_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5872_ _5998_/S _5872_/B vssd1 vssd1 vccd1 vccd1 _5872_/X sky130_fd_sc_hd__or2_1
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7611_ _7611_/CLK _7611_/D vssd1 vssd1 vccd1 vccd1 _7611_/Q sky130_fd_sc_hd__dfxtp_1
X_4823_ _4820_/X _7129_/Q _4835_/S vssd1 vssd1 vccd1 vccd1 _4824_/A sky130_fd_sc_hd__mux2_1
X_7542_ _7542_/CLK _7542_/D vssd1 vssd1 vccd1 vccd1 _7542_/Q sky130_fd_sc_hd__dfxtp_2
X_4754_ _4566_/X _7160_/Q _4760_/S vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__mux2_1
X_7473_ _7473_/CLK _7473_/D vssd1 vssd1 vccd1 vccd1 _7473_/Q sky130_fd_sc_hd__dfxtp_1
X_3705_ _3542_/X _7631_/Q _3707_/S vssd1 vssd1 vccd1 vccd1 _3706_/A sky130_fd_sc_hd__mux2_1
X_4685_ _4685_/A vssd1 vssd1 vccd1 vccd1 _7215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3636_ _3577_/A _3513_/A _3611_/A vssd1 vssd1 vccd1 vccd1 _6222_/A sky130_fd_sc_hd__a21oi_4
XFILLER_115_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3567_ _7354_/Q _7349_/Q vssd1 vssd1 vccd1 vccd1 _4376_/B sky130_fd_sc_hd__xnor2_1
XFILLER_115_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5306_ _5351_/A _5302_/X _5305_/X _5178_/X vssd1 vssd1 vccd1 vccd1 _5306_/X sky130_fd_sc_hd__o211a_1
Xclkbuf_0__3104_ _6401_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3104_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_88_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3498_ _7104_/Q vssd1 vssd1 vccd1 vccd1 _3511_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5237_ _5235_/X _5236_/X _5112_/X vssd1 vssd1 vccd1 vccd1 _5238_/B sky130_fd_sc_hd__o21ai_1
XFILLER_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5168_ _5257_/A _5168_/B vssd1 vssd1 vccd1 vccd1 _5168_/X sky130_fd_sc_hd__or2_1
X_5099_ _7202_/Q _5104_/B vssd1 vssd1 vccd1 vccd1 _5100_/A sky130_fd_sc_hd__and2_1
X_6436__67 _6438__69/A vssd1 vssd1 vccd1 vccd1 _7489_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4119_ _4118_/X _7448_/Q _4119_/S vssd1 vssd1 vccd1 vccd1 _4120_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4470_ _4473_/A _4473_/B vssd1 vssd1 vccd1 vccd1 _4474_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3075_ clkbuf_0__3075_/X vssd1 vssd1 vccd1 vccd1 _6357_/A sky130_fd_sc_hd__clkbuf_16
X_6140_ _6134_/Y _6135_/X _6775_/A _6775_/B vssd1 vssd1 vccd1 vccd1 _6157_/A sky130_fd_sc_hd__a211o_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5022_/A _5024_/B vssd1 vssd1 vccd1 vccd1 _5023_/A sky130_fd_sc_hd__and2_1
XFILLER_112_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6973_ _5440_/A _3501_/X _5380_/B _5587_/B _5586_/C vssd1 vssd1 vccd1 vccd1 _7010_/B
+ sky130_fd_sc_hd__a2111oi_4
X_5924_ _5924_/A vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5855_ _5855_/A vssd1 vssd1 vccd1 vccd1 _6005_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4806_ _4566_/X _7136_/Q _4812_/S vssd1 vssd1 vccd1 vccd1 _4807_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7516_/CLK sky130_fd_sc_hd__clkbuf_8
X_5786_ _7202_/Q _5029_/A _5794_/S vssd1 vssd1 vccd1 vccd1 _5787_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7525_ _7525_/CLK _7525_/D vssd1 vssd1 vccd1 vccd1 _7525_/Q sky130_fd_sc_hd__dfxtp_1
X_4737_ _4737_/A vssd1 vssd1 vccd1 vccd1 _7168_/D sky130_fd_sc_hd__clkbuf_1
X_4668_ _3807_/X _7230_/Q _4670_/S vssd1 vssd1 vccd1 vccd1 _4669_/A sky130_fd_sc_hd__mux2_1
X_7456_ _7456_/CLK _7456_/D vssd1 vssd1 vccd1 vccd1 _7456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6407_ _6413_/A vssd1 vssd1 vccd1 vccd1 _6407_/X sky130_fd_sc_hd__buf_1
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3619_ _3619_/A vssd1 vssd1 vccd1 vccd1 _7697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4599_ _4599_/A vssd1 vssd1 vccd1 vccd1 _7261_/D sky130_fd_sc_hd__clkbuf_1
X_7387_ _7387_/CLK _7387_/D vssd1 vssd1 vccd1 vccd1 _7387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5690__246 _5691__247/A vssd1 vssd1 vccd1 vccd1 _7140_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3281_ clkbuf_0__3281_/X vssd1 vssd1 vccd1 vccd1 _6698__137/A sky130_fd_sc_hd__clkbuf_16
XFILLER_13_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _3970_/A vssd1 vssd1 vccd1 vccd1 _7532_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__2713_ clkbuf_0__2713_/X vssd1 vssd1 vccd1 vccd1 _5687__244/A sky130_fd_sc_hd__clkbuf_16
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5640_ _7102_/Q _7201_/Q _6076_/S vssd1 vssd1 vccd1 vccd1 _5641_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5571_ _6579_/B _6610_/B _6569_/A _5570_/X vssd1 vssd1 vccd1 vccd1 _7071_/D sky130_fd_sc_hd__o211a_1
X_7310_ _7310_/CLK _7310_/D vssd1 vssd1 vccd1 vccd1 _7310_/Q sky130_fd_sc_hd__dfxtp_2
X_4522_ _7294_/Q _4343_/X _4522_/S vssd1 vssd1 vccd1 vccd1 _4523_/A sky130_fd_sc_hd__mux2_1
X_7241_ _7241_/CLK _7241_/D vssd1 vssd1 vccd1 vccd1 _7241_/Q sky130_fd_sc_hd__dfxtp_1
X_4453_ _3671_/A _4443_/B _4452_/Y vssd1 vssd1 vccd1 vccd1 _7315_/D sky130_fd_sc_hd__a21oi_1
X_7172_ _7172_/CLK _7172_/D vssd1 vssd1 vccd1 vccd1 _7172_/Q sky130_fd_sc_hd__dfxtp_1
X_4384_ _4384_/A _4391_/B vssd1 vssd1 vccd1 vccd1 _4388_/B sky130_fd_sc_hd__and2_1
XFILLER_86_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3058_ clkbuf_0__3058_/X vssd1 vssd1 vccd1 vccd1 _6210__386/A sky130_fd_sc_hd__clkbuf_16
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6446_/A vssd1 vssd1 vccd1 vccd1 _6452_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5005_/A vssd1 vssd1 vccd1 vccd1 _5005_/X sky130_fd_sc_hd__clkbuf_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6702__140 _6704__142/A vssd1 vssd1 vccd1 vccd1 _7584_/CLK sky130_fd_sc_hd__inv_2
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5907_ _5912_/A vssd1 vssd1 vccd1 vccd1 _5907_/X sky130_fd_sc_hd__clkbuf_4
X_6887_ _6170_/C _6879_/B _7658_/Q vssd1 vssd1 vccd1 vccd1 _6887_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5838_ _7582_/Q _7574_/Q _7566_/Q _7480_/Q _5870_/A _5857_/A vssd1 vssd1 vccd1 vccd1
+ _5838_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5769_ _5769_/A vssd1 vssd1 vccd1 vccd1 _7194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7508_ _7510_/CLK _7508_/D vssd1 vssd1 vccd1 vccd1 _7508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7439_ _7439_/CLK _7439_/D vssd1 vssd1 vccd1 vccd1 _7439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6321__455 _6323__457/A vssd1 vssd1 vccd1 vccd1 _7397_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6810_ _6859_/C vssd1 vssd1 vccd1 vccd1 _6868_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3953_ _3908_/X _7539_/Q _3957_/S vssd1 vssd1 vccd1 vccd1 _3954_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3884_ _3884_/A vssd1 vssd1 vccd1 vccd1 _7565_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__2627_ clkbuf_0__2627_/X vssd1 vssd1 vccd1 vccd1 _6972__4/A sky130_fd_sc_hd__clkbuf_16
XFILLER_31_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5623_ _5623_/A vssd1 vssd1 vccd1 vccd1 _7094_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3421_ _6957_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3421_/X sky130_fd_sc_hd__clkbuf_16
X_5554_ _7070_/Q _7069_/Q _6993_/A vssd1 vssd1 vccd1 vccd1 _5554_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5485_ _5481_/X _7203_/Q input20/X _5482_/X vssd1 vssd1 vccd1 vccd1 _5485_/X sky130_fd_sc_hd__a22o_2
X_4505_ _4505_/A vssd1 vssd1 vccd1 vccd1 _7302_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3283_ _6707_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3283_/X sky130_fd_sc_hd__clkbuf_16
X_4436_ _4436_/A vssd1 vssd1 vccd1 vccd1 _4443_/B sky130_fd_sc_hd__clkbuf_2
X_7224_ _7516_/CLK _7224_/D vssd1 vssd1 vccd1 vccd1 _7224_/Q sky130_fd_sc_hd__dfxtp_1
X_7155_ _7155_/CLK _7155_/D vssd1 vssd1 vccd1 vccd1 _7155_/Q sky130_fd_sc_hd__dfxtp_1
X_4367_ _7350_/Q vssd1 vssd1 vccd1 vccd1 _4368_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _7718_/Q _7653_/Q vssd1 vssd1 vccd1 vccd1 _6792_/B sky130_fd_sc_hd__xnor2_2
X_4298_ _4298_/A vssd1 vssd1 vccd1 vccd1 _7377_/D sky130_fd_sc_hd__clkbuf_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _7088_/CLK _7086_/D vssd1 vssd1 vccd1 vccd1 _7086_/Q sky130_fd_sc_hd__dfxtp_1
X_6037_ _6049_/A vssd1 vssd1 vccd1 vccd1 _6037_/X sky130_fd_sc_hd__buf_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6939_ _6951_/A vssd1 vssd1 vccd1 vccd1 _6939_/X sky130_fd_sc_hd__buf_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6953__41 _6956__44/A vssd1 vssd1 vccd1 vccd1 _7697_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6054__334 _6054__334/A vssd1 vssd1 vccd1 vccd1 _7260_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6709__146 _6712__149/A vssd1 vssd1 vccd1 vccd1 _7590_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6245__397 _6246__398/A vssd1 vssd1 vccd1 vccd1 _7337_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput106 _5094_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput139 _5032_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput128 _5009_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[15] sky130_fd_sc_hd__buf_2
Xoutput117 _5061_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[6] sky130_fd_sc_hd__buf_2
XFILLER_114_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5705__259 _5705__259/A vssd1 vssd1 vccd1 vccd1 _7153_/CLK sky130_fd_sc_hd__inv_2
X_5270_ _5270_/A vssd1 vssd1 vccd1 vccd1 _5290_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4221_ _4220_/X _7405_/Q _4227_/S vssd1 vssd1 vccd1 vccd1 _4222_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4152_ _4152_/A vssd1 vssd1 vccd1 vccd1 _7434_/D sky130_fd_sc_hd__clkbuf_1
X_4083_ _4083_/A vssd1 vssd1 vccd1 vccd1 _7461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6632__84 _6632__84/A vssd1 vssd1 vccd1 vccd1 _7528_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4985_ _4985_/A vssd1 vssd1 vccd1 vccd1 _4985_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3936_ _3936_/A vssd1 vssd1 vccd1 vccd1 _7547_/D sky130_fd_sc_hd__clkbuf_1
X_3867_ _3867_/A vssd1 vssd1 vccd1 vccd1 _7572_/D sky130_fd_sc_hd__clkbuf_1
X_3798_ _3820_/S vssd1 vssd1 vccd1 vccd1 _3811_/S sky130_fd_sc_hd__clkbuf_2
X_5606_ _5606_/A vssd1 vssd1 vccd1 vccd1 _7086_/D sky130_fd_sc_hd__clkbuf_1
X_6586_ _7509_/Q _6586_/B _6586_/C vssd1 vssd1 vccd1 vccd1 _6592_/B sky130_fd_sc_hd__and3_1
X_5537_ _5552_/S vssd1 vssd1 vccd1 vccd1 _5546_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_117_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5468_ _6463_/A _5438_/X _5449_/A _5467_/X vssd1 vssd1 vccd1 vccd1 _5468_/X sky130_fd_sc_hd__a31o_1
X_7207_ _7510_/CLK _7207_/D vssd1 vssd1 vccd1 vccd1 _7207_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3266_ _6619_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3266_/X sky130_fd_sc_hd__clkbuf_16
X_5399_ _5252_/X _5399_/B vssd1 vssd1 vccd1 vccd1 _5399_/X sky130_fd_sc_hd__and2b_1
X_4419_ _4434_/S vssd1 vssd1 vccd1 vccd1 _4428_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7138_ _7138_/CLK _7138_/D vssd1 vssd1 vccd1 vccd1 _7138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7069_ _7732_/CLK _7069_/D vssd1 vssd1 vccd1 vccd1 _7069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3101_ clkbuf_0__3101_/X vssd1 vssd1 vccd1 vccd1 _6413_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput19 caravel_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_2
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6681__124 _6681__124/A vssd1 vssd1 vccd1 vccd1 _7568_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__2961_ clkbuf_0__2961_/X vssd1 vssd1 vccd1 vccd1 _6067__344/A sky130_fd_sc_hd__clkbuf_16
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4770_ _7152_/Q _4325_/X _4774_/S vssd1 vssd1 vccd1 vccd1 _4771_/A sky130_fd_sc_hd__mux2_1
X_5711__263 _5711__263/A vssd1 vssd1 vccd1 vccd1 _7157_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ _3721_/A vssd1 vssd1 vccd1 vccd1 _7626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3652_ _4572_/A vssd1 vssd1 vccd1 vccd1 _3652_/X sky130_fd_sc_hd__clkbuf_2
X_3583_ _7706_/Q _3549_/X _3595_/S vssd1 vssd1 vccd1 vccd1 _3584_/A sky130_fd_sc_hd__mux2_1
X_5322_ _4384_/A _5315_/Y _5317_/Y _5319_/Y _5321_/Y vssd1 vssd1 vccd1 vccd1 _5322_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_88_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6334__465 _6337__468/A vssd1 vssd1 vccd1 vccd1 _7407_/CLK sky130_fd_sc_hd__inv_2
X_5253_ _7370_/Q _7341_/Q _7333_/Q _7296_/Q _4381_/A _5252_/X vssd1 vssd1 vccd1 vccd1
+ _5253_/X sky130_fd_sc_hd__mux4_2
X_4204_ _4204_/A vssd1 vssd1 vccd1 vccd1 _7411_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3051_ _6176_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3051_/X sky130_fd_sc_hd__clkbuf_16
X_5184_ _6274_/B vssd1 vssd1 vccd1 vccd1 _5184_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4135_ _4115_/X _7441_/Q _4137_/S vssd1 vssd1 vccd1 vccd1 _4136_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ _3911_/X _7468_/Q _4068_/S vssd1 vssd1 vccd1 vccd1 _4067_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4968_ _5092_/A vssd1 vssd1 vccd1 vccd1 _5106_/B sky130_fd_sc_hd__clkbuf_4
X_6707_ _6713_/A vssd1 vssd1 vccd1 vccd1 _6707_/X sky130_fd_sc_hd__buf_1
X_3919_ _3919_/A vssd1 vssd1 vccd1 vccd1 _7552_/D sky130_fd_sc_hd__clkbuf_1
X_7687_ _7687_/CLK _7687_/D vssd1 vssd1 vccd1 vccd1 _7687_/Q sky130_fd_sc_hd__dfxtp_1
X_4899_ _4899_/A vssd1 vssd1 vccd1 vccd1 _7072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6569_ _6569_/A vssd1 vssd1 vccd1 vccd1 _6569_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5654__217 _5655__218/A vssd1 vssd1 vccd1 vccd1 _7111_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3091_ clkbuf_0__3091_/X vssd1 vssd1 vccd1 vccd1 _6337__468/A sky130_fd_sc_hd__clkbuf_16
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5940_ _5938_/X _5939_/X _5998_/S vssd1 vssd1 vccd1 vccd1 _5940_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6067__344 _6067__344/A vssd1 vssd1 vccd1 vccd1 _7270_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5871_ _7393_/Q _7235_/Q _7551_/Q _7457_/Q _5857_/A _5870_/X vssd1 vssd1 vccd1 vccd1
+ _5872_/B sky130_fd_sc_hd__mux4_1
X_7610_ _7610_/CLK _7610_/D vssd1 vssd1 vccd1 vccd1 _7610_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4822_ _4844_/S vssd1 vssd1 vccd1 vccd1 _4835_/S sky130_fd_sc_hd__buf_2
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7541_ _7541_/CLK _7541_/D vssd1 vssd1 vccd1 vccd1 _7541_/Q sky130_fd_sc_hd__dfxtp_1
X_4753_ _4753_/A vssd1 vssd1 vccd1 vccd1 _7161_/D sky130_fd_sc_hd__clkbuf_1
X_7472_ _7472_/CLK _7472_/D vssd1 vssd1 vccd1 vccd1 _7472_/Q sky130_fd_sc_hd__dfxtp_1
X_3704_ _3704_/A vssd1 vssd1 vccd1 vccd1 _7632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4684_ _3804_/X _7215_/Q _4688_/S vssd1 vssd1 vccd1 vccd1 _4685_/A sky130_fd_sc_hd__mux2_1
X_3635_ _3983_/B _3926_/A _4301_/C vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__or3_4
XFILLER_108_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__3289_ clkbuf_0__3289_/X vssd1 vssd1 vccd1 vccd1 _6741__172/A sky130_fd_sc_hd__clkbuf_16
X_3566_ _7353_/Q _3570_/C vssd1 vssd1 vccd1 vccd1 _3756_/A sky130_fd_sc_hd__and2_1
XFILLER_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3497_ _7316_/Q vssd1 vssd1 vccd1 vccd1 _3822_/A sky130_fd_sc_hd__clkbuf_2
X_5305_ _5418_/A _5305_/B vssd1 vssd1 vccd1 vccd1 _5305_/X sky130_fd_sc_hd__or2_1
Xclkbuf_0__3103_ _6395_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3103_/X sky130_fd_sc_hd__clkbuf_16
X_5236_ _5236_/A vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5167_ _7526_/Q _7106_/Q _7558_/Q _7122_/Q _5132_/X _5135_/X vssd1 vssd1 vccd1 vccd1
+ _5168_/B sky130_fd_sc_hd__mux4_1
X_5098_ _5098_/A vssd1 vssd1 vccd1 vccd1 _5098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4118_ _7667_/Q vssd1 vssd1 vccd1 vccd1 _4118_/X sky130_fd_sc_hd__buf_2
X_4049_ _4049_/A vssd1 vssd1 vccd1 vccd1 _7476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5718__269 _5718__269/A vssd1 vssd1 vccd1 vccd1 _7163_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3074_ clkbuf_0__3074_/X vssd1 vssd1 vccd1 vccd1 _6259__409/A sky130_fd_sc_hd__clkbuf_16
XFILLER_97_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5021_/A vssd1 vssd1 vccd1 vccd1 _5021_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5923_ _5923_/A _5923_/B vssd1 vssd1 vccd1 vccd1 _5923_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6184__365 _6186__367/A vssd1 vssd1 vccd1 vccd1 _7295_/CLK sky130_fd_sc_hd__inv_2
X_6694__134 _6694__134/A vssd1 vssd1 vccd1 vccd1 _7578_/CLK sky130_fd_sc_hd__inv_2
X_5854_ _6003_/A _5854_/B vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__or2_1
X_6441__71 _6441__71/A vssd1 vssd1 vccd1 vccd1 _7493_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4805_ _4805_/A vssd1 vssd1 vccd1 vccd1 _7137_/D sky130_fd_sc_hd__clkbuf_1
X_7524_ _7524_/CLK _7524_/D vssd1 vssd1 vccd1 vccd1 _7524_/Q sky130_fd_sc_hd__dfxtp_2
X_5785_ _5800_/S vssd1 vssd1 vccd1 vccd1 _5794_/S sky130_fd_sc_hd__buf_2
X_4736_ _7168_/Q _4325_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4737_/A sky130_fd_sc_hd__mux2_1
X_4667_ _4667_/A vssd1 vssd1 vccd1 vccd1 _7231_/D sky130_fd_sc_hd__clkbuf_1
X_7455_ _7455_/CLK _7455_/D vssd1 vssd1 vccd1 vccd1 _7455_/Q sky130_fd_sc_hd__dfxtp_1
X_3618_ _3522_/X _7697_/Q _3624_/S vssd1 vssd1 vccd1 vccd1 _3619_/A sky130_fd_sc_hd__mux2_1
X_7386_ _7386_/CLK _7386_/D vssd1 vssd1 vccd1 vccd1 _7386_/Q sky130_fd_sc_hd__dfxtp_1
X_4598_ _4252_/X _7261_/Q _4598_/S vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3549_ _7328_/Q vssd1 vssd1 vccd1 vccd1 _3549_/X sky130_fd_sc_hd__clkbuf_8
X_6268_ _6277_/A vssd1 vssd1 vccd1 vccd1 _6268_/X sky130_fd_sc_hd__buf_1
X_5219_ _5319_/A _5219_/B vssd1 vssd1 vccd1 vccd1 _5219_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3280_ clkbuf_0__3280_/X vssd1 vssd1 vccd1 vccd1 _6691__131/A sky130_fd_sc_hd__clkbuf_16
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2712_ clkbuf_0__2712_/X vssd1 vssd1 vccd1 vccd1 _5679__237/A sky130_fd_sc_hd__clkbuf_16
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5570_ _7496_/Q _5570_/B _6609_/A vssd1 vssd1 vccd1 vccd1 _5570_/X sky130_fd_sc_hd__or3b_1
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4521_ _4521_/A vssd1 vssd1 vccd1 vccd1 _7295_/D sky130_fd_sc_hd__clkbuf_1
X_7240_ _7240_/CLK _7240_/D vssd1 vssd1 vccd1 vccd1 _7240_/Q sky130_fd_sc_hd__dfxtp_1
X_4452_ _3671_/A _4443_/B _4486_/C vssd1 vssd1 vccd1 vccd1 _4452_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7171_ _7171_/CLK _7171_/D vssd1 vssd1 vccd1 vccd1 _7171_/Q sky130_fd_sc_hd__dfxtp_1
X_4383_ _5315_/A _5331_/A _4393_/B vssd1 vssd1 vccd1 vccd1 _4391_/B sky130_fd_sc_hd__and3_1
XFILLER_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6122_ _6486_/B _6486_/C _6816_/A vssd1 vssd1 vccd1 vccd1 _6122_/X sky130_fd_sc_hd__a21o_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3057_ clkbuf_0__3057_/X vssd1 vssd1 vccd1 vccd1 _6254_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5004_/A _5012_/B vssd1 vssd1 vccd1 vccd1 _5005_/A sky130_fd_sc_hd__and2_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5906_ _7537_/Q _7678_/Q _7694_/Q _7280_/Q _5851_/X _5905_/X vssd1 vssd1 vccd1 vccd1
+ _5906_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6886_ _6886_/A vssd1 vssd1 vccd1 vccd1 _6886_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5837_ _7534_/Q _7675_/Q _7691_/Q _7277_/Q _5870_/A _5857_/A vssd1 vssd1 vccd1 vccd1
+ _5837_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5768_ _5010_/A _7194_/Q _5776_/S vssd1 vssd1 vccd1 vccd1 _5769_/A sky130_fd_sc_hd__mux2_1
X_4719_ _4719_/A vssd1 vssd1 vccd1 vccd1 _7176_/D sky130_fd_sc_hd__clkbuf_1
X_7507_ _7510_/CLK _7507_/D vssd1 vssd1 vccd1 vccd1 _7507_/Q sky130_fd_sc_hd__dfxtp_1
X_7438_ _7438_/CLK _7438_/D vssd1 vssd1 vccd1 vccd1 _7438_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7369_ _7369_/CLK _7369_/D vssd1 vssd1 vccd1 vccd1 _7369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3952_ _3952_/A vssd1 vssd1 vccd1 vccd1 _7540_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__2626_ clkbuf_0__2626_/X vssd1 vssd1 vccd1 vccd1 _5706_/A sky130_fd_sc_hd__clkbuf_16
X_3883_ _7565_/Q _3549_/X _3891_/S vssd1 vssd1 vccd1 vccd1 _3884_/A sky130_fd_sc_hd__mux2_1
X_5622_ _7094_/Q _7193_/Q _5624_/S vssd1 vssd1 vccd1 vccd1 _5623_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3420_ _6951_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3420_/X sky130_fd_sc_hd__clkbuf_16
X_5553_ _5553_/A vssd1 vssd1 vccd1 vccd1 _7068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4504_ _4235_/X _7302_/Q _4504_/S vssd1 vssd1 vccd1 vccd1 _4505_/A sky130_fd_sc_hd__mux2_1
X_5484_ _5481_/X _7202_/Q input19/X _5482_/X vssd1 vssd1 vccd1 vccd1 _5484_/X sky130_fd_sc_hd__a22o_2
Xclkbuf_0__3282_ _6701_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3282_/X sky130_fd_sc_hd__clkbuf_16
X_7223_ _7516_/CLK _7223_/D vssd1 vssd1 vccd1 vccd1 _7223_/Q sky130_fd_sc_hd__dfxtp_1
X_4435_ _4435_/A vssd1 vssd1 vccd1 vccd1 _7331_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__3109_ clkbuf_0__3109_/X vssd1 vssd1 vccd1 vccd1 _6426__59/A sky130_fd_sc_hd__clkbuf_16
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7154_ _7154_/CLK _7154_/D vssd1 vssd1 vccd1 vccd1 _7154_/Q sky130_fd_sc_hd__dfxtp_1
X_4366_ _7351_/Q vssd1 vssd1 vccd1 vccd1 _5337_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _6462_/A _6159_/A _6446_/B _6159_/C vssd1 vssd1 vccd1 vccd1 _6107_/A sky130_fd_sc_hd__or4_1
XFILLER_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4297_ _4258_/X _7377_/Q _4299_/S vssd1 vssd1 vccd1 vccd1 _4298_/A sky130_fd_sc_hd__mux2_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _7088_/CLK _7085_/D vssd1 vssd1 vccd1 vccd1 _7085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ _6938_/A vssd1 vssd1 vccd1 vccd1 _6938_/X sky130_fd_sc_hd__buf_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6869_ _6869_/A vssd1 vssd1 vccd1 vccd1 _7653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6061__339 _6061__339/A vssd1 vssd1 vccd1 vccd1 _7265_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput107 _5096_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput129 _5011_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[16] sky130_fd_sc_hd__buf_2
Xoutput118 _5063_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[7] sky130_fd_sc_hd__buf_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4220_ _4569_/A vssd1 vssd1 vccd1 vccd1 _4220_/X sky130_fd_sc_hd__buf_2
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ _7434_/Q _3597_/X _4155_/S vssd1 vssd1 vccd1 vccd1 _4152_/A sky130_fd_sc_hd__mux2_1
X_4082_ _7461_/Q _3804_/X _4086_/S vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6263__410 _6264__411/A vssd1 vssd1 vccd1 vccd1 _7350_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4984_ _6917_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4985_/A sky130_fd_sc_hd__and2_1
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3935_ _3648_/X _7547_/Q _3939_/S vssd1 vssd1 vccd1 vccd1 _3936_/A sky130_fd_sc_hd__mux2_1
X_3866_ _3735_/X _7572_/Q _3872_/S vssd1 vssd1 vccd1 vccd1 _3867_/A sky130_fd_sc_hd__mux2_1
X_5605_ _7086_/Q _5062_/A _5613_/S vssd1 vssd1 vccd1 vccd1 _5606_/A sky130_fd_sc_hd__mux2_1
X_3797_ _6236_/B _4606_/B _3797_/C vssd1 vssd1 vccd1 vccd1 _3820_/S sky130_fd_sc_hd__and3_4
X_6585_ _6583_/X _6584_/X _6569_/X vssd1 vssd1 vccd1 vccd1 _7508_/D sky130_fd_sc_hd__o21a_1
X_5536_ _5536_/A _5784_/B vssd1 vssd1 vccd1 vccd1 _5552_/S sky130_fd_sc_hd__nand2_2
XFILLER_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5467_ _5458_/X _7193_/Q input9/X _5102_/D vssd1 vssd1 vccd1 vccd1 _5467_/X sky130_fd_sc_hd__a22o_1
X_7206_ _7510_/CLK _7206_/D vssd1 vssd1 vccd1 vccd1 _7206_/Q sky130_fd_sc_hd__dfxtp_1
X_4418_ _4864_/A _4506_/B vssd1 vssd1 vccd1 vccd1 _4434_/S sky130_fd_sc_hd__or2_2
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5398_ _7523_/Q _7144_/Q _5429_/S vssd1 vssd1 vccd1 vccd1 _5399_/B sky130_fd_sc_hd__mux2_1
X_7137_ _7137_/CLK _7137_/D vssd1 vssd1 vccd1 vccd1 _7137_/Q sky130_fd_sc_hd__dfxtp_1
X_4349_ _7357_/Q _7358_/Q _4347_/Y _6220_/B vssd1 vssd1 vccd1 vccd1 _7357_/D sky130_fd_sc_hd__o211a_1
X_7068_ _7359_/CLK _7068_/D vssd1 vssd1 vccd1 vccd1 _7068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__3100_ clkbuf_0__3100_/X vssd1 vssd1 vccd1 vccd1 _6387__509/A sky130_fd_sc_hd__clkbuf_16
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6715__151 _6716__152/A vssd1 vssd1 vccd1 vccd1 _7595_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2960_ clkbuf_0__2960_/X vssd1 vssd1 vccd1 vccd1 _6060__338/A sky130_fd_sc_hd__clkbuf_16
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3720_ _3530_/X _7626_/Q _3722_/S vssd1 vssd1 vccd1 vccd1 _3721_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3651_ _7325_/Q vssd1 vssd1 vccd1 vccd1 _4572_/A sky130_fd_sc_hd__clkbuf_4
X_3582_ _3604_/S vssd1 vssd1 vccd1 vccd1 _3595_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6370_ _6370_/A vssd1 vssd1 vccd1 vccd1 _6370_/X sky130_fd_sc_hd__buf_1
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5321_ _5315_/A _5320_/X _4384_/A vssd1 vssd1 vccd1 vccd1 _5321_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5252_ _5252_/A vssd1 vssd1 vccd1 vccd1 _5252_/X sky130_fd_sc_hd__clkbuf_4
X_4203_ _4109_/X _7411_/Q _4203_/S vssd1 vssd1 vccd1 vccd1 _4204_/A sky130_fd_sc_hd__mux2_1
X_5183_ _5187_/A _5380_/B _5183_/C _5587_/C vssd1 vssd1 vccd1 vccd1 _6274_/B sky130_fd_sc_hd__or4_2
XFILLER_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4134_ _4134_/A vssd1 vssd1 vccd1 vccd1 _7442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4065_ _4065_/A vssd1 vssd1 vccd1 vccd1 _7469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _4967_/A vssd1 vssd1 vccd1 vccd1 _4967_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3918_ _3917_/X _7552_/Q _3924_/S vssd1 vssd1 vccd1 vccd1 _3919_/A sky130_fd_sc_hd__mux2_1
X_7686_ _7686_/CLK _7686_/D vssd1 vssd1 vccd1 vccd1 _7686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4898_ _4843_/X _7072_/Q _4898_/S vssd1 vssd1 vccd1 vccd1 _4899_/A sky130_fd_sc_hd__mux2_1
X_3849_ _3849_/A vssd1 vssd1 vccd1 vccd1 _7579_/D sky130_fd_sc_hd__clkbuf_1
X_6568_ _7505_/Q _6589_/B _6594_/C vssd1 vssd1 vccd1 vccd1 _6568_/X sky130_fd_sc_hd__and3_1
XFILLER_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6499_ _6567_/A vssd1 vssd1 vccd1 vccd1 _6579_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__3090_ clkbuf_0__3090_/X vssd1 vssd1 vccd1 vccd1 _6332__464/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5870_ _5870_/A vssd1 vssd1 vccd1 vccd1 _5870_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4821_ _4821_/A _4864_/B vssd1 vssd1 vccd1 vccd1 _4844_/S sky130_fd_sc_hd__or2_2
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7540_ _7540_/CLK _7540_/D vssd1 vssd1 vccd1 vccd1 _7540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4752_ _4560_/X _7161_/Q _4760_/S vssd1 vssd1 vccd1 vccd1 _4753_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7471_ _7471_/CLK _7471_/D vssd1 vssd1 vccd1 vccd1 _7471_/Q sky130_fd_sc_hd__dfxtp_1
X_4683_ _4683_/A vssd1 vssd1 vccd1 vccd1 _7216_/D sky130_fd_sc_hd__clkbuf_1
X_3703_ _3538_/X _7632_/Q _3707_/S vssd1 vssd1 vccd1 vccd1 _3704_/A sky130_fd_sc_hd__mux2_1
X_6340__470 _6342__472/A vssd1 vssd1 vccd1 vccd1 _7412_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3634_ _4561_/B vssd1 vssd1 vccd1 vccd1 _4301_/C sky130_fd_sc_hd__clkinv_2
Xclkbuf_1_0__f__3288_ clkbuf_0__3288_/X vssd1 vssd1 vccd1 vccd1 _6737__169/A sky130_fd_sc_hd__clkbuf_16
X_3565_ _3565_/A vssd1 vssd1 vccd1 vccd1 _5230_/B sky130_fd_sc_hd__inv_2
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3496_ _3609_/A vssd1 vssd1 vccd1 vccd1 _4436_/A sky130_fd_sc_hd__clkbuf_2
X_5304_ _7371_/Q _7342_/Q _7334_/Q _7297_/Q _5403_/S _5303_/X vssd1 vssd1 vccd1 vccd1
+ _5305_/B sky130_fd_sc_hd__mux4_1
Xclkbuf_0__3102_ _6389_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3102_/X sky130_fd_sc_hd__clkbuf_16
X_5235_ _6487_/A vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_102_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5166_ _5418_/A vssd1 vssd1 vccd1 vccd1 _5257_/A sky130_fd_sc_hd__clkbuf_2
X_5097_ _7201_/Q _5104_/B vssd1 vssd1 vccd1 vccd1 _5098_/A sky130_fd_sc_hd__and2_1
X_4117_ _4117_/A vssd1 vssd1 vccd1 vccd1 _7449_/D sky130_fd_sc_hd__clkbuf_1
X_4048_ _3911_/X _7476_/Q _4050_/S vssd1 vssd1 vccd1 vccd1 _4049_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _5995_/X _5998_/X _5999_/S vssd1 vssd1 vccd1 vccd1 _5999_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7669_ _7674_/CLK _7669_/D vssd1 vssd1 vccd1 vccd1 _7669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5660__222 _5661__223/A vssd1 vssd1 vccd1 vccd1 _7116_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__3073_ clkbuf_0__3073_/X vssd1 vssd1 vccd1 vccd1 _6252__403/A sky130_fd_sc_hd__clkbuf_16
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5020_/A _5024_/B vssd1 vssd1 vccd1 vccd1 _5021_/A sky130_fd_sc_hd__and2_1
XFILLER_85_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6728__161 _6729__162/A vssd1 vssd1 vccd1 vccd1 _7605_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5922_ _7395_/Q _7237_/Q _7553_/Q _7459_/Q _5921_/X _4468_/A vssd1 vssd1 vccd1 vccd1
+ _5923_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5853_ _7583_/Q _7575_/Q _7567_/Q _7481_/Q _5851_/X _5852_/X vssd1 vssd1 vccd1 vccd1
+ _5854_/B sky130_fd_sc_hd__mux4_2
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4804_ _4560_/X _7137_/Q _4812_/S vssd1 vssd1 vccd1 vccd1 _4805_/A sky130_fd_sc_hd__mux2_1
X_5784_ _5784_/A _5784_/B vssd1 vssd1 vccd1 vccd1 _5800_/S sky130_fd_sc_hd__and2_4
X_7523_ _7523_/CLK _7523_/D vssd1 vssd1 vccd1 vccd1 _7523_/Q sky130_fd_sc_hd__dfxtp_2
X_4735_ _4735_/A vssd1 vssd1 vccd1 vccd1 _7169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4666_ _3804_/X _7231_/Q _4670_/S vssd1 vssd1 vccd1 vccd1 _4667_/A sky130_fd_sc_hd__mux2_1
X_7454_ _7454_/CLK _7454_/D vssd1 vssd1 vccd1 vccd1 _7454_/Q sky130_fd_sc_hd__dfxtp_1
X_4597_ _4597_/A vssd1 vssd1 vccd1 vccd1 _7262_/D sky130_fd_sc_hd__clkbuf_1
X_3617_ _3617_/A vssd1 vssd1 vccd1 vccd1 _7698_/D sky130_fd_sc_hd__clkbuf_1
X_7385_ _7385_/CLK _7385_/D vssd1 vssd1 vccd1 vccd1 _7385_/Q sky130_fd_sc_hd__dfxtp_1
X_3548_ _3548_/A vssd1 vssd1 vccd1 vccd1 _7707_/D sky130_fd_sc_hd__clkbuf_1
X_5724__274 _5724__274/A vssd1 vssd1 vccd1 vccd1 _7168_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3479_ _7317_/Q _7312_/Q vssd1 vssd1 vccd1 vccd1 _3484_/B sky130_fd_sc_hd__xor2_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5218_ _7287_/Q _7073_/Q _7700_/Q _7361_/Q _5173_/A _5171_/X vssd1 vssd1 vccd1 vccd1
+ _5219_/B sky130_fd_sc_hd__mux4_1
XFILLER_96_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5149_ _7368_/Q _7339_/Q _7331_/Q _7294_/Q _5397_/S _5148_/X vssd1 vssd1 vccd1 vccd1
+ _5150_/B sky130_fd_sc_hd__mux4_1
XFILLER_72_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6347__476 _6347__476/A vssd1 vssd1 vccd1 vccd1 _7418_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6250__401 _6253__404/A vssd1 vssd1 vccd1 vccd1 _7341_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5521__192 _5523__194/A vssd1 vssd1 vccd1 vccd1 _7049_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2711_ clkbuf_0__2711_/X vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_63_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5667__228 _5667__228/A vssd1 vssd1 vccd1 vccd1 _7122_/CLK sky130_fd_sc_hd__inv_2
X_4520_ _7295_/Q _4340_/X _4522_/S vssd1 vssd1 vccd1 vccd1 _4521_/A sky130_fd_sc_hd__mux2_1
X_4451_ _4451_/A vssd1 vssd1 vccd1 vccd1 _7316_/D sky130_fd_sc_hd__clkbuf_1
X_7170_ _7170_/CLK _7170_/D vssd1 vssd1 vccd1 vccd1 _7170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__3056_ clkbuf_0__3056_/X vssd1 vssd1 vccd1 vccd1 _6204__382/A sky130_fd_sc_hd__clkbuf_16
X_6121_ _6816_/A _6486_/B _6486_/C vssd1 vssd1 vccd1 vccd1 _6121_/Y sky130_fd_sc_hd__nand3_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4382_ _5381_/A _7359_/Q _4382_/C vssd1 vssd1 vccd1 vccd1 _4393_/B sky130_fd_sc_hd__and3b_1
XFILLER_98_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6190__370 _6191__371/A vssd1 vssd1 vccd1 vccd1 _7300_/CLK sky130_fd_sc_hd__inv_2
X_5003_ _5106_/B vssd1 vssd1 vccd1 vccd1 _5012_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5905_ _5908_/A vssd1 vssd1 vccd1 vccd1 _5905_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6965__51 _6968__54/A vssd1 vssd1 vccd1 vccd1 _7707_/CLK sky130_fd_sc_hd__inv_2
X_6885_ _6885_/A vssd1 vssd1 vccd1 vccd1 _7657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5836_ _5921_/A vssd1 vssd1 vccd1 vccd1 _5857_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5767_ _5782_/S vssd1 vssd1 vccd1 vccd1 _5776_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4718_ _4566_/X _7176_/Q _4724_/S vssd1 vssd1 vccd1 vccd1 _4719_/A sky130_fd_sc_hd__mux2_1
X_7506_ _7510_/CLK _7506_/D vssd1 vssd1 vccd1 vccd1 _7506_/Q sky130_fd_sc_hd__dfxtp_1
X_4649_ _4649_/A vssd1 vssd1 vccd1 vccd1 _7239_/D sky130_fd_sc_hd__clkbuf_1
X_7437_ _7437_/CLK _7437_/D vssd1 vssd1 vccd1 vccd1 _7437_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7368_ _7368_/CLK _7368_/D vssd1 vssd1 vccd1 vccd1 _7368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7299_ _7299_/CLK _7299_/D vssd1 vssd1 vccd1 vccd1 _7299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6644__94 _6644__94/A vssd1 vssd1 vccd1 vccd1 _7538_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3951_ _3905_/X _7540_/Q _3957_/S vssd1 vssd1 vccd1 vccd1 _3952_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2625_ clkbuf_0__2625_/X vssd1 vssd1 vccd1 vccd1 _6938_/A sky130_fd_sc_hd__clkbuf_16
X_6670_ _6682_/A vssd1 vssd1 vccd1 vccd1 _6670_/X sky130_fd_sc_hd__buf_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3882_ _3897_/S vssd1 vssd1 vccd1 vccd1 _3891_/S sky130_fd_sc_hd__clkbuf_2
X_5621_ _5621_/A vssd1 vssd1 vccd1 vccd1 _7093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5552_ _6923_/A _7068_/Q _5552_/S vssd1 vssd1 vccd1 vccd1 _5553_/A sky130_fd_sc_hd__mux2_1
X_4503_ _4503_/A vssd1 vssd1 vccd1 vccd1 _7303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6257__407 _6259__409/A vssd1 vssd1 vccd1 vccd1 _7347_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5483_ _5481_/X _7201_/Q input18/X _5482_/X vssd1 vssd1 vccd1 vccd1 _5483_/X sky130_fd_sc_hd__a22o_2
Xclkbuf_0__3281_ _6695_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3281_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7222_ _7516_/CLK _7222_/D vssd1 vssd1 vccd1 vccd1 _7222_/Q sky130_fd_sc_hd__dfxtp_1
X_4434_ _4235_/X _7331_/Q _4434_/S vssd1 vssd1 vccd1 vccd1 _4435_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3108_ clkbuf_0__3108_/X vssd1 vssd1 vccd1 vccd1 _6619_/A sky130_fd_sc_hd__clkbuf_16
X_5528__198 _5528__198/A vssd1 vssd1 vccd1 vccd1 _7055_/CLK sky130_fd_sc_hd__inv_2
X_7153_ _7153_/CLK _7153_/D vssd1 vssd1 vccd1 vccd1 _7153_/Q sky130_fd_sc_hd__dfxtp_1
X_4365_ _4365_/A vssd1 vssd1 vccd1 vccd1 _7352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7084_ _7088_/CLK _7084_/D vssd1 vssd1 vccd1 vccd1 _7084_/Q sky130_fd_sc_hd__dfxtp_1
X_6104_ _7723_/Q _7722_/Q _7721_/Q _7720_/Q vssd1 vssd1 vccd1 vccd1 _6159_/C sky130_fd_sc_hd__or4_4
XFILLER_100_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4296_ _4296_/A vssd1 vssd1 vccd1 vccd1 _7378_/D sky130_fd_sc_hd__clkbuf_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6868_ _6868_/A _6868_/B _6868_/C vssd1 vssd1 vccd1 vccd1 _6869_/A sky130_fd_sc_hd__and3_1
X_5819_ _5924_/A vssd1 vssd1 vccd1 vccd1 _5819_/X sky130_fd_sc_hd__buf_4
X_6799_ _6889_/B _6780_/Y _6795_/Y _6798_/X vssd1 vssd1 vccd1 vccd1 _7638_/D sky130_fd_sc_hd__o211a_1
XFILLER_6_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6197__376 _6200__379/A vssd1 vssd1 vccd1 vccd1 _7306_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6403__521 _6403__521/A vssd1 vssd1 vccd1 vccd1 _7463_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput108 _5098_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput119 _5065_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[8] sky130_fd_sc_hd__buf_2
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4150_ _4150_/A vssd1 vssd1 vccd1 vccd1 _7435_/D sky130_fd_sc_hd__clkbuf_1
X_4081_ _4081_/A vssd1 vssd1 vccd1 vccd1 _7462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4983_ _4983_/A vssd1 vssd1 vccd1 vccd1 _4983_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3934_ _3934_/A vssd1 vssd1 vccd1 vccd1 _7548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3865_ _3865_/A vssd1 vssd1 vccd1 vccd1 _7573_/D sky130_fd_sc_hd__clkbuf_1
X_6304__441 _6304__441/A vssd1 vssd1 vccd1 vccd1 _7383_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5604_ _5637_/A vssd1 vssd1 vccd1 vccd1 _5613_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_118_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3796_ _3822_/A _3861_/C _3796_/C vssd1 vssd1 vccd1 vccd1 _4606_/B sky130_fd_sc_hd__and3_2
X_6584_ _6586_/B _6589_/B _6594_/C vssd1 vssd1 vccd1 vccd1 _6584_/X sky130_fd_sc_hd__and3_1
XFILLER_11_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5535_ _7070_/Q _5535_/B _7069_/Q vssd1 vssd1 vccd1 vccd1 _5784_/B sky130_fd_sc_hd__nor3b_4
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5466_ _7717_/Q vssd1 vssd1 vccd1 vccd1 _6463_/A sky130_fd_sc_hd__clkbuf_4
X_7205_ _7516_/CLK _7205_/D vssd1 vssd1 vccd1 vccd1 _7205_/Q sky130_fd_sc_hd__dfxtp_2
X_4417_ _4417_/A vssd1 vssd1 vccd1 vccd1 _7339_/D sky130_fd_sc_hd__clkbuf_1
X_5397_ _7160_/Q _7152_/Q _5397_/S vssd1 vssd1 vccd1 vccd1 _5397_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7136_ _7136_/CLK _7136_/D vssd1 vssd1 vccd1 vccd1 _7136_/Q sky130_fd_sc_hd__dfxtp_1
X_4348_ _6222_/A vssd1 vssd1 vccd1 vccd1 _6220_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4279_ _7385_/Q _3600_/X _4281_/S vssd1 vssd1 vccd1 vccd1 _4280_/A sky130_fd_sc_hd__mux2_1
X_7067_ _7359_/CLK _7067_/D vssd1 vssd1 vccd1 vccd1 _7067_/Q sky130_fd_sc_hd__dfxtp_1
X_6018_ _6018_/A vssd1 vssd1 vccd1 vccd1 _6018_/X sky130_fd_sc_hd__buf_1
XFILLER_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6205__383 _6206__384/A vssd1 vssd1 vccd1 vccd1 _7313_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6722__156 _6725__159/A vssd1 vssd1 vccd1 vccd1 _7600_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3650_ _3650_/A vssd1 vssd1 vccd1 vccd1 _7688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3581_ _4882_/A _4400_/A vssd1 vssd1 vccd1 vccd1 _3604_/S sky130_fd_sc_hd__nor2_2
XFILLER_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5320_ _7174_/Q _7306_/Q _7492_/Q _7182_/Q _5148_/X _4382_/C vssd1 vssd1 vccd1 vccd1
+ _5320_/X sky130_fd_sc_hd__mux4_1
X_5251_ _7348_/Q vssd1 vssd1 vccd1 vccd1 _5252_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4202_ _4202_/A vssd1 vssd1 vccd1 vccd1 _7412_/D sky130_fd_sc_hd__clkbuf_1
X_5182_ _7084_/Q _7083_/Q vssd1 vssd1 vccd1 vccd1 _5587_/C sky130_fd_sc_hd__or2b_1
XFILLER_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4133_ _4112_/X _7442_/Q _4137_/S vssd1 vssd1 vccd1 vccd1 _4134_/A sky130_fd_sc_hd__mux2_1
X_4064_ _3908_/X _7469_/Q _4068_/S vssd1 vssd1 vccd1 vccd1 _4065_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4966_ _5748_/A _4966_/B vssd1 vssd1 vccd1 vccd1 _4967_/A sky130_fd_sc_hd__and2_1
X_3917_ _3917_/A vssd1 vssd1 vccd1 vccd1 _3917_/X sky130_fd_sc_hd__buf_4
X_7685_ _7685_/CLK _7685_/D vssd1 vssd1 vccd1 vccd1 _7685_/Q sky130_fd_sc_hd__dfxtp_1
X_4897_ _4897_/A vssd1 vssd1 vccd1 vccd1 _7073_/D sky130_fd_sc_hd__clkbuf_1
X_3848_ _3738_/X _7579_/Q _3852_/S vssd1 vssd1 vccd1 vccd1 _3849_/A sky130_fd_sc_hd__mux2_1
X_3779_ _3779_/A vssd1 vssd1 vccd1 vccd1 _7605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6567_ _6567_/A vssd1 vssd1 vccd1 vccd1 _6594_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5518_ _5518_/A vssd1 vssd1 vccd1 vccd1 _5518_/X sky130_fd_sc_hd__buf_1
Xclkbuf_4_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7359_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_105_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6498_ _6498_/A vssd1 vssd1 vccd1 vccd1 _6567_/A sky130_fd_sc_hd__clkbuf_2
X_5449_ _5449_/A vssd1 vssd1 vccd1 vccd1 _5449_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7119_ _7119_/CLK _7119_/D vssd1 vssd1 vccd1 vccd1 _7119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4820_ _7328_/Q vssd1 vssd1 vccd1 vccd1 _4820_/X sky130_fd_sc_hd__buf_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4766_/S vssd1 vssd1 vccd1 vccd1 _4760_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_119_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7470_ _7470_/CLK _7470_/D vssd1 vssd1 vccd1 vccd1 _7470_/Q sky130_fd_sc_hd__dfxtp_1
X_4682_ _3801_/X _7216_/Q _4688_/S vssd1 vssd1 vccd1 vccd1 _4683_/A sky130_fd_sc_hd__mux2_1
X_3702_ _3702_/A vssd1 vssd1 vccd1 vccd1 _7633_/D sky130_fd_sc_hd__clkbuf_1
X_6421_ _6427_/A vssd1 vssd1 vccd1 vccd1 _6421_/X sky130_fd_sc_hd__buf_1
X_3633_ _4560_/A vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3287_ clkbuf_0__3287_/X vssd1 vssd1 vccd1 vccd1 _6731__164/A sky130_fd_sc_hd__clkbuf_16
X_3564_ _4350_/A _4376_/C vssd1 vssd1 vccd1 vccd1 _3565_/A sky130_fd_sc_hd__xor2_1
X_5303_ _5303_/A vssd1 vssd1 vccd1 vccd1 _5303_/X sky130_fd_sc_hd__clkbuf_4
X_3495_ _5584_/B _7329_/Q vssd1 vssd1 vccd1 vccd1 _3609_/A sky130_fd_sc_hd__and2b_1
X_6283_ _6289_/A vssd1 vssd1 vccd1 vccd1 _6283_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3101_ _6388_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3101_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_69_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5234_ _7731_/Q vssd1 vssd1 vccd1 vccd1 _6487_/A sky130_fd_sc_hd__clkbuf_2
X_5165_ _5351_/A _5165_/B vssd1 vssd1 vccd1 vccd1 _5165_/X sky130_fd_sc_hd__or2_1
X_4116_ _4115_/X _7449_/Q _4119_/S vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5096_ _5096_/A vssd1 vssd1 vccd1 vccd1 _5096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4047_ _4047_/A vssd1 vssd1 vccd1 vccd1 _7477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5996_/X _5997_/X _5998_/S vssd1 vssd1 vccd1 vccd1 _5998_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4949_ _4949_/A vssd1 vssd1 vccd1 vccd1 _7038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7668_ _7670_/CLK _7668_/D vssd1 vssd1 vccd1 vccd1 _7668_/Q sky130_fd_sc_hd__dfxtp_2
X_6619_ _6619_/A vssd1 vssd1 vccd1 vccd1 _6619_/X sky130_fd_sc_hd__buf_1
XFILLER_20_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7599_ _7599_/CLK _7599_/D vssd1 vssd1 vccd1 vccd1 _7599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__3072_ clkbuf_0__3072_/X vssd1 vssd1 vccd1 vccd1 _6247__399/A sky130_fd_sc_hd__clkbuf_16
XFILLER_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5921_ _5921_/A vssd1 vssd1 vccd1 vccd1 _5921_/X sky130_fd_sc_hd__buf_2
XFILLER_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5852_ _5908_/A vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__buf_4
X_4803_ _4818_/S vssd1 vssd1 vccd1 vccd1 _4812_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5783_ _5783_/A vssd1 vssd1 vccd1 vccd1 _7201_/D sky130_fd_sc_hd__clkbuf_1
X_7522_ _7522_/CLK _7522_/D vssd1 vssd1 vccd1 vccd1 _7522_/Q sky130_fd_sc_hd__dfxtp_1
X_4734_ _7169_/Q _4320_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4735_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4665_ _4665_/A vssd1 vssd1 vccd1 vccd1 _7232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7453_ _7453_/CLK _7453_/D vssd1 vssd1 vccd1 vccd1 _7453_/Q sky130_fd_sc_hd__dfxtp_1
X_4596_ _4249_/X _7262_/Q _4598_/S vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__mux2_1
X_3616_ _3469_/X _7698_/Q _3624_/S vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__mux2_1
X_7384_ _7384_/CLK _7384_/D vssd1 vssd1 vccd1 vccd1 _7384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3547_ _3546_/X _7707_/Q _3547_/S vssd1 vssd1 vccd1 vccd1 _3548_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3478_ _7316_/Q _3822_/C vssd1 vssd1 vccd1 vccd1 _3484_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5217_ _5433_/A _5217_/B _5217_/C vssd1 vssd1 vccd1 vccd1 _5217_/Y sky130_fd_sc_hd__nor3_1
XFILLER_56_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5148_ _5148_/A vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__buf_2
XFILLER_28_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5079_ _7193_/Q _5079_/B vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__and2_1
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2710_ clkbuf_0__2710_/X vssd1 vssd1 vccd1 vccd1 _5673__233/A sky130_fd_sc_hd__clkbuf_16
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4450_ _4606_/B _4450_/B _4486_/C vssd1 vssd1 vccd1 vccd1 _4451_/A sky130_fd_sc_hd__and3b_1
X_4381_ _4381_/A vssd1 vssd1 vccd1 vccd1 _4382_/C sky130_fd_sc_hd__buf_2
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3055_ clkbuf_0__3055_/X vssd1 vssd1 vccd1 vccd1 _6200__379/A sky130_fd_sc_hd__clkbuf_16
X_6120_ _5235_/X _6119_/B _5281_/X vssd1 vssd1 vccd1 vccd1 _6486_/C sky130_fd_sc_hd__o21ai_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/A vssd1 vssd1 vccd1 vccd1 _5002_/X sky130_fd_sc_hd__clkbuf_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5904_ _7220_/Q _5814_/X _5903_/Y _5880_/X vssd1 vssd1 vccd1 vccd1 _7220_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6884_ _6886_/A _6884_/B _6884_/C vssd1 vssd1 vccd1 vccd1 _6885_/A sky130_fd_sc_hd__and3_1
XFILLER_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5835_ _5912_/A vssd1 vssd1 vccd1 vccd1 _5870_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5766_ _5766_/A _5784_/B vssd1 vssd1 vccd1 vccd1 _5782_/S sky130_fd_sc_hd__nand2_4
XFILLER_108_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4717_ _4717_/A vssd1 vssd1 vccd1 vccd1 _7177_/D sky130_fd_sc_hd__clkbuf_1
X_7505_ _7510_/CLK _7505_/D vssd1 vssd1 vccd1 vccd1 _7505_/Q sky130_fd_sc_hd__dfxtp_1
X_4648_ _4246_/X _7239_/Q _4652_/S vssd1 vssd1 vccd1 vccd1 _4649_/A sky130_fd_sc_hd__mux2_1
X_7436_ _7436_/CLK _7436_/D vssd1 vssd1 vccd1 vccd1 _7436_/Q sky130_fd_sc_hd__dfxtp_1
X_4579_ _4578_/X _7268_/Q _4585_/S vssd1 vssd1 vccd1 vccd1 _4580_/A sky130_fd_sc_hd__mux2_1
X_7367_ _7367_/CLK _7367_/D vssd1 vssd1 vccd1 vccd1 _7367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6353__481 _6356__484/A vssd1 vssd1 vccd1 vccd1 _7423_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7298_ _7298_/CLK _7298_/D vssd1 vssd1 vccd1 vccd1 _7298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6677__120 _6681__124/A vssd1 vssd1 vccd1 vccd1 _7564_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_14_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7510_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_75_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5673__233 _5673__233/A vssd1 vssd1 vccd1 vccd1 _7127_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3950_ _3950_/A vssd1 vssd1 vccd1 vccd1 _7541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3881_ _4400_/A _4864_/B vssd1 vssd1 vccd1 vccd1 _3897_/S sky130_fd_sc_hd__nor2_4
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5620_ _7093_/Q _5077_/A _5624_/S vssd1 vssd1 vccd1 vccd1 _5621_/A sky130_fd_sc_hd__mux2_1
X_5551_ _5551_/A vssd1 vssd1 vccd1 vccd1 _7067_/D sky130_fd_sc_hd__clkbuf_1
X_4502_ _4232_/X _7303_/Q _4504_/S vssd1 vssd1 vccd1 vccd1 _4503_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7221_ _7516_/CLK _7221_/D vssd1 vssd1 vccd1 vccd1 _7221_/Q sky130_fd_sc_hd__dfxtp_1
X_5482_ _5482_/A vssd1 vssd1 vccd1 vccd1 _5482_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3280_ _6689_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3280_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f__3107_ clkbuf_0__3107_/X vssd1 vssd1 vccd1 vccd1 _6719_/A sky130_fd_sc_hd__clkbuf_16
X_4433_ _4433_/A vssd1 vssd1 vccd1 vccd1 _7332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7152_ _7152_/CLK _7152_/D vssd1 vssd1 vccd1 vccd1 _7152_/Q sky130_fd_sc_hd__dfxtp_1
X_4364_ _4364_/A _6272_/C _4364_/C vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__and3_1
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4295_ _4255_/X _7378_/Q _4299_/S vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7083_ _7088_/CLK _7083_/D vssd1 vssd1 vccd1 vccd1 _7083_/Q sky130_fd_sc_hd__dfxtp_1
X_6103_ _6127_/C vssd1 vssd1 vccd1 vccd1 _6446_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6867_ _7653_/Q _6870_/C vssd1 vssd1 vccd1 vccd1 _6868_/C sky130_fd_sc_hd__nand2_1
X_5818_ _5912_/A vssd1 vssd1 vccd1 vccd1 _5818_/X sky130_fd_sc_hd__buf_6
X_6798_ _6800_/A _6794_/A _6781_/X _6886_/A vssd1 vssd1 vccd1 vccd1 _6798_/X sky130_fd_sc_hd__o31a_1
X_5749_ _5764_/S vssd1 vssd1 vccd1 vccd1 _5758_/S sky130_fd_sc_hd__clkbuf_2
X_7419_ _7419_/CLK _7419_/D vssd1 vssd1 vccd1 vccd1 _7419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput109 _5100_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[24] sky130_fd_sc_hd__buf_2
XFILLER_114_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5744__289 _5744__289/A vssd1 vssd1 vccd1 vccd1 _7183_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4080_ _7462_/Q _3801_/X _4086_/S vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__2959_ clkbuf_0__2959_/X vssd1 vssd1 vccd1 vccd1 _6056_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4982_ _6915_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4983_/A sky130_fd_sc_hd__and2_1
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3933_ _3644_/X _7548_/Q _3939_/S vssd1 vssd1 vccd1 vccd1 _3934_/A sky130_fd_sc_hd__mux2_1
X_3864_ _3730_/X _7573_/Q _3872_/S vssd1 vssd1 vccd1 vccd1 _3865_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5603_ _5603_/A vssd1 vssd1 vccd1 vccd1 _7085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3795_ _4606_/A vssd1 vssd1 vccd1 vccd1 _6236_/B sky130_fd_sc_hd__buf_2
X_6583_ _6587_/B _6583_/B _6583_/C vssd1 vssd1 vccd1 vccd1 _6583_/X sky130_fd_sc_hd__and3b_1
XCaravelHost_230 vssd1 vssd1 vccd1 vccd1 core1Index[0] CaravelHost_230/LO sky130_fd_sc_hd__conb_1
X_5465_ _7718_/Q _5438_/X _5449_/A _5464_/X vssd1 vssd1 vccd1 vccd1 _5465_/X sky130_fd_sc_hd__a31o_1
XFILLER_105_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7204_ _7516_/CLK _7204_/D vssd1 vssd1 vccd1 vccd1 _7204_/Q sky130_fd_sc_hd__dfxtp_2
X_6270__416 _6275__418/A vssd1 vssd1 vccd1 vccd1 _7356_/CLK sky130_fd_sc_hd__inv_2
X_4416_ _7339_/Q _4343_/X _4416_/S vssd1 vssd1 vccd1 vccd1 _4417_/A sky130_fd_sc_hd__mux2_1
X_7135_ _7135_/CLK _7135_/D vssd1 vssd1 vccd1 vccd1 _7135_/Q sky130_fd_sc_hd__dfxtp_1
X_5396_ _5396_/A _5396_/B vssd1 vssd1 vccd1 vccd1 _5396_/X sky130_fd_sc_hd__or2_1
XFILLER_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4347_ _4350_/B vssd1 vssd1 vccd1 vccd1 _4347_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4278_ _4278_/A vssd1 vssd1 vccd1 vccd1 _7386_/D sky130_fd_sc_hd__clkbuf_1
X_7066_ _7359_/CLK _7066_/D vssd1 vssd1 vccd1 vccd1 _7066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6919_ _6919_/A _6923_/B vssd1 vssd1 vccd1 vccd1 _6920_/A sky130_fd_sc_hd__and2_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5808__297 _5808__297/A vssd1 vssd1 vccd1 vccd1 _7215_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6212__388 _6213__389/A vssd1 vssd1 vccd1 vccd1 _7318_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6366__491 _6369__494/A vssd1 vssd1 vccd1 vccd1 _7433_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3580_ _4918_/A vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__3089_ clkbuf_0__3089_/X vssd1 vssd1 vccd1 vccd1 _6351_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5250_ _5351_/A _5250_/B vssd1 vssd1 vccd1 vccd1 _5250_/Y sky130_fd_sc_hd__nor2_1
X_4201_ _4106_/X _7412_/Q _4203_/S vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5181_ _5131_/X _5165_/X _5168_/X _5179_/X _5433_/A vssd1 vssd1 vccd1 vccd1 _5181_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_96_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4132_ _4132_/A vssd1 vssd1 vccd1 vccd1 _7443_/D sky130_fd_sc_hd__clkbuf_1
X_4063_ _4063_/A vssd1 vssd1 vccd1 vccd1 _7470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4965_ _4965_/A vssd1 vssd1 vccd1 vccd1 _4965_/X sky130_fd_sc_hd__clkbuf_1
X_6766__17 _6766__17/A vssd1 vssd1 vccd1 vccd1 _7636_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3916_ _3916_/A vssd1 vssd1 vccd1 vccd1 _7553_/D sky130_fd_sc_hd__clkbuf_1
X_6083__352 _6083__352/A vssd1 vssd1 vccd1 vccd1 _7281_/CLK sky130_fd_sc_hd__inv_2
X_6044__325 _6046__327/A vssd1 vssd1 vccd1 vccd1 _7251_/CLK sky130_fd_sc_hd__inv_2
X_7684_ _7684_/CLK _7684_/D vssd1 vssd1 vccd1 vccd1 _7684_/Q sky130_fd_sc_hd__dfxtp_1
X_5686__243 _5686__243/A vssd1 vssd1 vccd1 vccd1 _7137_/CLK sky130_fd_sc_hd__inv_2
X_4896_ _4840_/X _7073_/Q _4898_/S vssd1 vssd1 vccd1 vccd1 _4897_/A sky130_fd_sc_hd__mux2_1
X_3847_ _3847_/A vssd1 vssd1 vccd1 vccd1 _7580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ _3730_/X _7605_/Q _3786_/S vssd1 vssd1 vccd1 vccd1 _3779_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6566_ _6566_/A _6566_/B _6571_/B vssd1 vssd1 vccd1 vccd1 _6566_/X sky130_fd_sc_hd__and3_1
X_6497_ _7496_/Q _6572_/A _6572_/B _6572_/C vssd1 vssd1 vccd1 vccd1 _6498_/A sky130_fd_sc_hd__and4_1
XFILLER_105_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5448_ _5494_/S vssd1 vssd1 vccd1 vccd1 _5448_/X sky130_fd_sc_hd__clkbuf_2
X_5379_ _5469_/A _7010_/A _5440_/A vssd1 vssd1 vccd1 vccd1 _5436_/B sky130_fd_sc_hd__and3_1
XFILLER_113_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7118_ _7118_/CLK _7118_/D vssd1 vssd1 vccd1 vccd1 _7118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7049_ _7049_/CLK _7049_/D vssd1 vssd1 vccd1 vccd1 _7049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4864_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _4766_/S sky130_fd_sc_hd__or2_2
X_4681_ _4681_/A vssd1 vssd1 vccd1 vccd1 _7217_/D sky130_fd_sc_hd__clkbuf_1
X_3701_ _3534_/X _7633_/Q _3701_/S vssd1 vssd1 vccd1 vccd1 _3702_/A sky130_fd_sc_hd__mux2_1
X_6420_ _6688_/A vssd1 vssd1 vccd1 vccd1 _6420_/X sky130_fd_sc_hd__buf_1
X_3632_ _7328_/Q vssd1 vssd1 vccd1 vccd1 _4560_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__3286_ clkbuf_0__3286_/X vssd1 vssd1 vccd1 vccd1 _6725__159/A sky130_fd_sc_hd__clkbuf_16
X_6351_ _6351_/A vssd1 vssd1 vccd1 vccd1 _6351_/X sky130_fd_sc_hd__buf_1
X_6416__532 _6416__532/A vssd1 vssd1 vccd1 vccd1 _7474_/CLK sky130_fd_sc_hd__inv_2
X_5302_ _7289_/Q _7075_/Q _7702_/Q _7363_/Q _5207_/X _5225_/X vssd1 vssd1 vccd1 vccd1
+ _5302_/X sky130_fd_sc_hd__mux4_1
X_3563_ _7356_/Q _7351_/Q vssd1 vssd1 vccd1 vccd1 _4376_/C sky130_fd_sc_hd__xnor2_1
X_3494_ _3494_/A _3494_/B _3494_/C _3494_/D vssd1 vssd1 vccd1 vccd1 _5584_/B sky130_fd_sc_hd__and4_4
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3100_ _6382_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3100_/X sky130_fd_sc_hd__clkbuf_16
X_5233_ _5217_/Y _5228_/X _5308_/A _5231_/X _5236_/A vssd1 vssd1 vccd1 vccd1 _5238_/A
+ sky130_fd_sc_hd__o311a_1
X_5164_ _7114_/Q _7162_/Q _7683_/Q _7606_/Q _5138_/X _5148_/X vssd1 vssd1 vccd1 vccd1
+ _5165_/B sky130_fd_sc_hd__mux4_1
XFILLER_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4115_ _7668_/Q vssd1 vssd1 vccd1 vccd1 _4115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5095_ _7200_/Q _5104_/B vssd1 vssd1 vccd1 vccd1 _5096_/A sky130_fd_sc_hd__and2_1
XFILLER_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4046_ _3908_/X _7477_/Q _4050_/S vssd1 vssd1 vccd1 vccd1 _4047_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _7249_/Q _7233_/Q _7479_/Q _7471_/Q _5860_/X _5870_/X vssd1 vssd1 vccd1 vccd1
+ _5997_/X sky130_fd_sc_hd__mux4_1
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4948_ _3813_/X _7038_/Q _4952_/S vssd1 vssd1 vccd1 vccd1 _4949_/A sky130_fd_sc_hd__mux2_1
X_6671__115 _6674__118/A vssd1 vssd1 vccd1 vccd1 _7559_/CLK sky130_fd_sc_hd__inv_2
X_7667_ _7674_/CLK _7667_/D vssd1 vssd1 vccd1 vccd1 _7667_/Q sky130_fd_sc_hd__dfxtp_1
X_4879_ _4879_/A vssd1 vssd1 vccd1 vccd1 _7107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7598_ _7598_/CLK _7598_/D vssd1 vssd1 vccd1 vccd1 _7598_/Q sky130_fd_sc_hd__dfxtp_1
X_6549_ _6553_/B _6553_/C vssd1 vssd1 vccd1 vccd1 _6550_/C sky130_fd_sc_hd__nand2_1
X_6317__452 _6317__452/A vssd1 vssd1 vccd1 vccd1 _7394_/CLK sky130_fd_sc_hd__inv_2
X_5508__186 _5509__187/A vssd1 vssd1 vccd1 vccd1 _7042_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5920_ _6005_/A _5920_/B vssd1 vssd1 vccd1 vccd1 _5920_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5533__202 _5572__204/A vssd1 vssd1 vccd1 vccd1 _7059_/CLK sky130_fd_sc_hd__inv_2
X_5851_ _5912_/A vssd1 vssd1 vccd1 vccd1 _5851_/X sky130_fd_sc_hd__clkbuf_8
X_4802_ _4802_/A _4918_/B vssd1 vssd1 vccd1 vccd1 _4818_/S sky130_fd_sc_hd__or2_2
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5782_ _5027_/A _7201_/Q _5782_/S vssd1 vssd1 vccd1 vccd1 _5783_/A sky130_fd_sc_hd__mux2_1
X_7521_ _7521_/CLK _7521_/D vssd1 vssd1 vccd1 vccd1 _7521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4733_ _4748_/S vssd1 vssd1 vccd1 vccd1 _4742_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_119_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6735__167 _6736__168/A vssd1 vssd1 vccd1 vccd1 _7611_/CLK sky130_fd_sc_hd__inv_2
X_7452_ _7452_/CLK _7452_/D vssd1 vssd1 vccd1 vccd1 _7452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4664_ _3801_/X _7232_/Q _4670_/S vssd1 vssd1 vccd1 vccd1 _4665_/A sky130_fd_sc_hd__mux2_1
X_4595_ _4595_/A vssd1 vssd1 vccd1 vccd1 _7263_/D sky130_fd_sc_hd__clkbuf_1
X_3615_ _3630_/S vssd1 vssd1 vccd1 vccd1 _3624_/S sky130_fd_sc_hd__clkbuf_2
X_7383_ _7383_/CLK _7383_/D vssd1 vssd1 vccd1 vccd1 _7383_/Q sky130_fd_sc_hd__dfxtp_1
X_3546_ _3923_/A vssd1 vssd1 vccd1 vccd1 _3546_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f__3269_ clkbuf_0__3269_/X vssd1 vssd1 vccd1 vccd1 _6638__89/A sky130_fd_sc_hd__clkbuf_16
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3477_ _7317_/Q _7316_/Q _7315_/Q vssd1 vssd1 vccd1 vccd1 _4443_/A sky130_fd_sc_hd__and3_1
X_5216_ _5209_/X _5214_/X _5215_/X _5289_/A _5158_/X vssd1 vssd1 vccd1 vccd1 _5217_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5147_ _5403_/S vssd1 vssd1 vccd1 vccd1 _5397_/S sky130_fd_sc_hd__buf_2
X_5078_ _5078_/A vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__clkbuf_1
X_4029_ _3911_/X _7484_/Q _4031_/S vssd1 vssd1 vccd1 vccd1 _4030_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7719_ _7722_/CLK _7719_/D vssd1 vssd1 vccd1 vccd1 _7719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6057__335 _6061__339/A vssd1 vssd1 vccd1 vccd1 _7261_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4380_ _5421_/S vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__3054_ clkbuf_0__3054_/X vssd1 vssd1 vccd1 vccd1 _6191__371/A sky130_fd_sc_hd__clkbuf_16
XFILLER_98_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5001_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _5002_/A sky130_fd_sc_hd__and2_1
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5903_ _5882_/X _5893_/X _5902_/Y _5814_/A vssd1 vssd1 vccd1 vccd1 _5903_/Y sky130_fd_sc_hd__o211ai_4
X_6883_ _6170_/C _6889_/B _6879_/B _6879_/C vssd1 vssd1 vccd1 vccd1 _6884_/C sky130_fd_sc_hd__o211ai_1
X_5834_ _7314_/Q vssd1 vssd1 vccd1 vccd1 _5902_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5765_ _5765_/A vssd1 vssd1 vccd1 vccd1 _7193_/D sky130_fd_sc_hd__clkbuf_1
X_4716_ _4560_/X _7177_/Q _4724_/S vssd1 vssd1 vccd1 vccd1 _4717_/A sky130_fd_sc_hd__mux2_1
X_7504_ _7652_/CLK _7504_/D vssd1 vssd1 vccd1 vccd1 _7504_/Q sky130_fd_sc_hd__dfxtp_1
X_4647_ _4647_/A vssd1 vssd1 vccd1 vccd1 _7240_/D sky130_fd_sc_hd__clkbuf_1
X_7435_ _7435_/CLK _7435_/D vssd1 vssd1 vccd1 vccd1 _7435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7366_ _7366_/CLK _7366_/D vssd1 vssd1 vccd1 vccd1 _7366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4578_ _4578_/A vssd1 vssd1 vccd1 vccd1 _4578_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3529_ _7671_/Q vssd1 vssd1 vccd1 vccd1 _3911_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7297_ _7297_/CLK _7297_/D vssd1 vssd1 vccd1 vccd1 _7297_/Q sky130_fd_sc_hd__dfxtp_1
X_6248_ _6254_/A vssd1 vssd1 vccd1 vccd1 _6248_/X sky130_fd_sc_hd__buf_1
XFILLER_57_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6360__486 _6360__486/A vssd1 vssd1 vccd1 vccd1 _7428_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3880_ _3983_/B _3926_/A _4561_/B vssd1 vssd1 vccd1 vccd1 _4864_/B sky130_fd_sc_hd__or3_4
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5550_ _6921_/A _7067_/Q _5552_/S vssd1 vssd1 vccd1 vccd1 _5551_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4501_ _4501_/A vssd1 vssd1 vccd1 vccd1 _7304_/D sky130_fd_sc_hd__clkbuf_1
X_5481_ _5481_/A vssd1 vssd1 vccd1 vccd1 _5481_/X sky130_fd_sc_hd__clkbuf_2
X_5680__238 _5681__239/A vssd1 vssd1 vccd1 vccd1 _7132_/CLK sky130_fd_sc_hd__inv_2
X_7220_ _7516_/CLK _7220_/D vssd1 vssd1 vccd1 vccd1 _7220_/Q sky130_fd_sc_hd__dfxtp_1
X_4432_ _4232_/X _7332_/Q _4434_/S vssd1 vssd1 vccd1 vccd1 _4433_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__3106_ clkbuf_0__3106_/X vssd1 vssd1 vccd1 vccd1 _6416__532/A sky130_fd_sc_hd__clkbuf_16
X_7151_ _7151_/CLK _7151_/D vssd1 vssd1 vccd1 vccd1 _7151_/Q sky130_fd_sc_hd__dfxtp_1
X_4363_ _4363_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _4364_/C sky130_fd_sc_hd__or2_1
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4294_ _4294_/A vssd1 vssd1 vccd1 vccd1 _7379_/D sky130_fd_sc_hd__clkbuf_1
X_7082_ _7088_/CLK _7082_/D vssd1 vssd1 vccd1 vccd1 _7082_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6127_/B vssd1 vssd1 vccd1 vccd1 _6159_/A sky130_fd_sc_hd__buf_2
XFILLER_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6650__99 _6650__99/A vssd1 vssd1 vccd1 vccd1 _7543_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6866_ _7653_/Q _6870_/C vssd1 vssd1 vccd1 vccd1 _6868_/B sky130_fd_sc_hd__or2_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5817_ _7310_/Q vssd1 vssd1 vccd1 vccd1 _5912_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6797_ _6797_/A vssd1 vssd1 vccd1 vccd1 _6886_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5748_ _5748_/A _5784_/B vssd1 vssd1 vccd1 vccd1 _5764_/S sky130_fd_sc_hd__nand2_2
X_7418_ _7418_/CLK _7418_/D vssd1 vssd1 vccd1 vccd1 _7418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7349_ _7349_/CLK _7349_/D vssd1 vssd1 vccd1 vccd1 _7349_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_104_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6944__34 _6944__34/A vssd1 vssd1 vccd1 vccd1 _7690_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6410__527 _6410__527/A vssd1 vssd1 vccd1 vccd1 _7469_/CLK sky130_fd_sc_hd__inv_2
Xoutput92 _7071_/Q vssd1 vssd1 vccd1 vccd1 caravel_uart_tx sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__2958_ clkbuf_0__2958_/X vssd1 vssd1 vccd1 vccd1 _6052__332/A sky130_fd_sc_hd__clkbuf_16
XFILLER_95_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _5106_/B vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6720_ _6744_/A vssd1 vssd1 vccd1 vccd1 _6720_/X sky130_fd_sc_hd__buf_1
X_3932_ _3932_/A vssd1 vssd1 vccd1 vccd1 _7549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3863_ _3878_/S vssd1 vssd1 vccd1 vccd1 _3872_/S sky130_fd_sc_hd__clkbuf_2
X_6651_ _6651_/A vssd1 vssd1 vccd1 vccd1 _6651_/X sky130_fd_sc_hd__buf_1
XFILLER_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5602_ _7085_/Q _5060_/A _5602_/S vssd1 vssd1 vccd1 vccd1 _5603_/A sky130_fd_sc_hd__mux2_1
X_6582_ _6586_/B _6586_/C vssd1 vssd1 vccd1 vccd1 _6583_/B sky130_fd_sc_hd__or2_1
X_3794_ _7674_/Q vssd1 vssd1 vccd1 vccd1 _3794_/X sky130_fd_sc_hd__buf_6
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XCaravelHost_220 vssd1 vssd1 vccd1 vccd1 CaravelHost_220/HI partID[3] sky130_fd_sc_hd__conb_1
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XCaravelHost_231 vssd1 vssd1 vccd1 vccd1 partID[0] CaravelHost_231/LO sky130_fd_sc_hd__conb_1
X_5464_ _5458_/X _7192_/Q _5102_/D input8/X vssd1 vssd1 vccd1 vccd1 _5464_/X sky130_fd_sc_hd__a22o_1
X_5395_ _7176_/Q _7308_/Q _7494_/Q _7184_/Q _5148_/A _5330_/S vssd1 vssd1 vccd1 vccd1
+ _5396_/B sky130_fd_sc_hd__mux4_1
X_7203_ _7525_/CLK _7203_/D vssd1 vssd1 vccd1 vccd1 _7203_/Q sky130_fd_sc_hd__dfxtp_1
X_4415_ _4415_/A vssd1 vssd1 vccd1 vccd1 _7340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7134_ _7134_/CLK _7134_/D vssd1 vssd1 vccd1 vccd1 _7134_/Q sky130_fd_sc_hd__dfxtp_1
X_4346_ _4363_/B vssd1 vssd1 vccd1 vccd1 _4350_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6311__447 _6312__448/A vssd1 vssd1 vccd1 vccd1 _7389_/CLK sky130_fd_sc_hd__inv_2
X_4277_ _7386_/Q _3597_/X _4281_/S vssd1 vssd1 vccd1 vccd1 _4278_/A sky130_fd_sc_hd__mux2_1
X_7065_ _7088_/CLK _7065_/D vssd1 vssd1 vccd1 vccd1 _7065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6918_ _6918_/A vssd1 vssd1 vccd1 vccd1 _7671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6849_ _7649_/Q _6849_/B vssd1 vssd1 vccd1 vccd1 _6850_/B sky130_fd_sc_hd__or2_1
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3088_ clkbuf_0__3088_/X vssd1 vssd1 vccd1 vccd1 _6323__457/A sky130_fd_sc_hd__clkbuf_16
XFILLER_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ _4200_/A vssd1 vssd1 vccd1 vccd1 _7413_/D sky130_fd_sc_hd__clkbuf_1
X_5180_ _7351_/Q vssd1 vssd1 vccd1 vccd1 _5433_/A sky130_fd_sc_hd__buf_2
XFILLER_110_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4131_ _4109_/X _7443_/Q _4131_/S vssd1 vssd1 vccd1 vccd1 _4132_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4062_ _3905_/X _7470_/Q _4068_/S vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5501__181 _5502__182/A vssd1 vssd1 vccd1 vccd1 _7037_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4964_ _5536_/A _4966_/B vssd1 vssd1 vccd1 vccd1 _4965_/A sky130_fd_sc_hd__and2_1
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3915_ _3914_/X _7553_/Q _3915_/S vssd1 vssd1 vccd1 vccd1 _3916_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7683_ _7683_/CLK _7683_/D vssd1 vssd1 vccd1 vccd1 _7683_/Q sky130_fd_sc_hd__dfxtp_2
X_4895_ _4895_/A vssd1 vssd1 vccd1 vccd1 _7074_/D sky130_fd_sc_hd__clkbuf_1
X_3846_ _3735_/X _7580_/Q _3852_/S vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3777_ _3792_/S vssd1 vssd1 vccd1 vccd1 _3786_/S sky130_fd_sc_hd__buf_2
X_6565_ _7505_/Q _6576_/D vssd1 vssd1 vccd1 vccd1 _6571_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6496_ _6594_/A _6503_/B _6466_/Y _6475_/X _6495_/X vssd1 vssd1 vccd1 vccd1 _6572_/C
+ sky130_fd_sc_hd__a2111oi_1
X_5447_ _7723_/Q vssd1 vssd1 vccd1 vccd1 _6137_/A sky130_fd_sc_hd__buf_4
X_5378_ _5592_/D vssd1 vssd1 vccd1 vccd1 _5469_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7117_ _7117_/CLK _7117_/D vssd1 vssd1 vccd1 vccd1 _7117_/Q sky130_fd_sc_hd__dfxtp_1
X_4329_ _7365_/Q _4328_/X _4335_/S vssd1 vssd1 vccd1 vccd1 _4330_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7048_ _7048_/CLK _7048_/D vssd1 vssd1 vccd1 vccd1 _7048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__2726_ clkbuf_0__2726_/X vssd1 vssd1 vccd1 vccd1 _5804__294/A sky130_fd_sc_hd__clkbuf_16
XFILLER_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _3700_/A vssd1 vssd1 vccd1 vccd1 _7634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ _3794_/X _7217_/Q _4688_/S vssd1 vssd1 vccd1 vccd1 _4681_/A sky130_fd_sc_hd__mux2_1
X_3631_ _3631_/A vssd1 vssd1 vccd1 vccd1 _7691_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__3285_ clkbuf_0__3285_/X vssd1 vssd1 vccd1 vccd1 _6732_/A sky130_fd_sc_hd__clkbuf_16
X_3562_ _7355_/Q _7354_/Q _7353_/Q _7352_/Q vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__and4_1
X_5301_ _5298_/X _5300_/X _5413_/A vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__mux2_1
X_3493_ _3493_/A _3493_/B vssd1 vssd1 vccd1 vccd1 _3494_/D sky130_fd_sc_hd__nor2_1
X_5232_ _5232_/A _5232_/B vssd1 vssd1 vccd1 vccd1 _5236_/A sky130_fd_sc_hd__or2_2
XFILLER_102_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5163_ _5163_/A vssd1 vssd1 vccd1 vccd1 _5351_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4114_ _4114_/A vssd1 vssd1 vccd1 vccd1 _7450_/D sky130_fd_sc_hd__clkbuf_1
X_5094_ _5094_/A vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__clkbuf_1
X_6050__330 _6052__332/A vssd1 vssd1 vccd1 vccd1 _7256_/CLK sky130_fd_sc_hd__inv_2
X_4045_ _4045_/A vssd1 vssd1 vccd1 vccd1 _7478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _7217_/Q _7043_/Q _7265_/Q _7257_/Q _5841_/X _5913_/X vssd1 vssd1 vccd1 vccd1
+ _5996_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4947_ _4947_/A vssd1 vssd1 vccd1 vccd1 _7039_/D sky130_fd_sc_hd__clkbuf_1
X_4878_ _4840_/X _7107_/Q _4880_/S vssd1 vssd1 vccd1 vccd1 _4879_/A sky130_fd_sc_hd__mux2_1
X_7666_ _7727_/CLK _7666_/D vssd1 vssd1 vccd1 vccd1 _7666_/Q sky130_fd_sc_hd__dfxtp_1
X_3829_ _3829_/A vssd1 vssd1 vccd1 vccd1 _7588_/D sky130_fd_sc_hd__clkbuf_1
X_6617_ _6515_/A _6615_/B _6615_/A vssd1 vssd1 vccd1 vccd1 _7516_/D sky130_fd_sc_hd__a21boi_1
X_7597_ _7597_/CLK _7597_/D vssd1 vssd1 vccd1 vccd1 _7597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6548_ _6553_/B _6553_/C vssd1 vssd1 vccd1 vccd1 _6550_/B sky130_fd_sc_hd__or2_1
XFILLER_118_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6479_ _6507_/B _6507_/C _6562_/A vssd1 vssd1 vccd1 vccd1 _6479_/X sky130_fd_sc_hd__a21bo_1
XINSDIODE2_0 _3920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5701__255 _5702__256/A vssd1 vssd1 vccd1 vccd1 _7149_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2709_ clkbuf_0__2709_/X vssd1 vssd1 vccd1 vccd1 _5667__228/A sky130_fd_sc_hd__clkbuf_16
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5850_ _5869_/A vssd1 vssd1 vccd1 vccd1 _6003_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4801_ _4801_/A vssd1 vssd1 vccd1 vccd1 _7138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5781_ _5781_/A vssd1 vssd1 vccd1 vccd1 _7200_/D sky130_fd_sc_hd__clkbuf_1
X_7520_ _7520_/CLK _7520_/D vssd1 vssd1 vccd1 vccd1 _7520_/Q sky130_fd_sc_hd__dfxtp_1
X_4732_ _4918_/A _4846_/A vssd1 vssd1 vccd1 vccd1 _4748_/S sky130_fd_sc_hd__nor2_2
X_4663_ _4663_/A vssd1 vssd1 vccd1 vccd1 _7233_/D sky130_fd_sc_hd__clkbuf_1
X_7451_ _7451_/CLK _7451_/D vssd1 vssd1 vccd1 vccd1 _7451_/Q sky130_fd_sc_hd__dfxtp_1
X_3614_ _4542_/B _4660_/A vssd1 vssd1 vccd1 vccd1 _3630_/S sky130_fd_sc_hd__nand2_2
X_4594_ _4246_/X _7263_/Q _4598_/S vssd1 vssd1 vccd1 vccd1 _4595_/A sky130_fd_sc_hd__mux2_1
X_7382_ _7382_/CLK _7382_/D vssd1 vssd1 vccd1 vccd1 _7382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3545_ _7667_/Q vssd1 vssd1 vccd1 vccd1 _3923_/A sky130_fd_sc_hd__buf_4
Xclkbuf_1_0__f__3268_ clkbuf_0__3268_/X vssd1 vssd1 vccd1 vccd1 _6632__84/A sky130_fd_sc_hd__clkbuf_16
X_6333_ _6333_/A vssd1 vssd1 vccd1 vccd1 _6333_/X sky130_fd_sc_hd__buf_1
XFILLER_115_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3476_ _3861_/C vssd1 vssd1 vccd1 vccd1 _3671_/A sky130_fd_sc_hd__clkbuf_2
X_5215_ _7171_/Q _7303_/Q _7489_/Q _7179_/Q _5173_/A _5171_/X vssd1 vssd1 vccd1 vccd1
+ _5215_/X sky130_fd_sc_hd__mux4_1
X_6195_ _6195_/A vssd1 vssd1 vccd1 vccd1 _6195_/X sky130_fd_sc_hd__buf_1
XFILLER_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5146_ _5245_/A vssd1 vssd1 vccd1 vccd1 _5403_/S sky130_fd_sc_hd__buf_2
X_5077_ _5077_/A _5079_/B vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__and2_1
X_4028_ _4028_/A vssd1 vssd1 vccd1 vccd1 _7485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6432__64 _6432__64/A vssd1 vssd1 vccd1 vccd1 _7486_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5979_ _5975_/X _5978_/X _5999_/S vssd1 vssd1 vccd1 vccd1 _5979_/X sky130_fd_sc_hd__mux2_2
XFILLER_100_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7718_ _7722_/CLK _7718_/D vssd1 vssd1 vccd1 vccd1 _7718_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7649_ _7655_/CLK _7649_/D vssd1 vssd1 vccd1 vccd1 _7649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5699__254 _5699__254/A vssd1 vssd1 vccd1 vccd1 _7148_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__3053_ clkbuf_0__3053_/X vssd1 vssd1 vccd1 vccd1 _6188__369/A sky130_fd_sc_hd__clkbuf_16
XFILLER_112_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5000_/A vssd1 vssd1 vccd1 vccd1 _5000_/X sky130_fd_sc_hd__clkbuf_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6741__172 _6741__172/A vssd1 vssd1 vccd1 vccd1 _7616_/CLK sky130_fd_sc_hd__inv_2
X_6951_ _6951_/A vssd1 vssd1 vccd1 vccd1 _6951_/X sky130_fd_sc_hd__buf_1
X_5902_ _5902_/A _5902_/B vssd1 vssd1 vccd1 vccd1 _5902_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6882_ _7656_/Q _6879_/B _7657_/Q vssd1 vssd1 vccd1 vccd1 _6884_/B sky130_fd_sc_hd__a21o_1
X_5833_ _5833_/A vssd1 vssd1 vccd1 vccd1 _5833_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5764_ _5008_/A _7193_/Q _5764_/S vssd1 vssd1 vccd1 vccd1 _5765_/A sky130_fd_sc_hd__mux2_1
X_7503_ _7652_/CLK _7503_/D vssd1 vssd1 vccd1 vccd1 _7503_/Q sky130_fd_sc_hd__dfxtp_1
X_4715_ _4730_/S vssd1 vssd1 vccd1 vccd1 _4724_/S sky130_fd_sc_hd__clkbuf_2
X_4646_ _4243_/X _7240_/Q _4652_/S vssd1 vssd1 vccd1 vccd1 _4647_/A sky130_fd_sc_hd__mux2_1
X_7434_ _7434_/CLK _7434_/D vssd1 vssd1 vccd1 vccd1 _7434_/Q sky130_fd_sc_hd__dfxtp_1
X_4577_ _4577_/A vssd1 vssd1 vccd1 vccd1 _7269_/D sky130_fd_sc_hd__clkbuf_1
X_7365_ _7365_/CLK _7365_/D vssd1 vssd1 vccd1 vccd1 _7365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3528_ _3528_/A vssd1 vssd1 vccd1 vccd1 _7712_/D sky130_fd_sc_hd__clkbuf_1
X_7296_ _7296_/CLK _7296_/D vssd1 vssd1 vccd1 vccd1 _7296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5129_ _5381_/A _5441_/D vssd1 vssd1 vccd1 vccd1 _5129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6063__340 _6065__342/A vssd1 vssd1 vccd1 vccd1 _7266_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6684__126 _6685__127/A vssd1 vssd1 vccd1 vccd1 _7570_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6752__5 _6756__9/A vssd1 vssd1 vccd1 vccd1 _7624_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5714__265 _5718__269/A vssd1 vssd1 vccd1 vccd1 _7159_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4500_ _4229_/X _7304_/Q _4504_/S vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5480_ _5474_/X _7200_/Q input17/X _5475_/X vssd1 vssd1 vccd1 vccd1 _5480_/X sky130_fd_sc_hd__a22o_2
X_4431_ _4431_/A vssd1 vssd1 vccd1 vccd1 _7333_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__3105_ clkbuf_0__3105_/X vssd1 vssd1 vccd1 vccd1 _6410__527/A sky130_fd_sc_hd__clkbuf_16
X_7150_ _7150_/CLK _7150_/D vssd1 vssd1 vccd1 vccd1 _7150_/Q sky130_fd_sc_hd__dfxtp_1
X_4362_ _4362_/A vssd1 vssd1 vccd1 vccd1 _7353_/D sky130_fd_sc_hd__clkbuf_1
X_4293_ _4252_/X _7379_/Q _4293_/S vssd1 vssd1 vccd1 vccd1 _4294_/A sky130_fd_sc_hd__mux2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7081_ _7088_/CLK _7081_/D vssd1 vssd1 vccd1 vccd1 _7081_/Q sky130_fd_sc_hd__dfxtp_2
X_6101_ _6163_/A _6492_/C _7650_/Q vssd1 vssd1 vccd1 vccd1 _6101_/X sky130_fd_sc_hd__a21bo_1
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6635__86 _6637__88/A vssd1 vssd1 vccd1 vccd1 _7530_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6865_ _7652_/Q _6857_/X _6864_/X vssd1 vssd1 vccd1 vccd1 _7652_/D sky130_fd_sc_hd__o21ba_1
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5816_ _5855_/A vssd1 vssd1 vccd1 vccd1 _5959_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_50_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6796_ input1/X vssd1 vssd1 vccd1 vccd1 _6800_/A sky130_fd_sc_hd__inv_2
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7417_ _7417_/CLK _7417_/D vssd1 vssd1 vccd1 vccd1 _7417_/Q sky130_fd_sc_hd__dfxtp_1
X_4629_ _4629_/A vssd1 vssd1 vccd1 vccd1 _7248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7348_ _7348_/CLK _7348_/D vssd1 vssd1 vccd1 vccd1 _7348_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7279_ _7279_/CLK _7279_/D vssd1 vssd1 vccd1 vccd1 _7279_/Q sky130_fd_sc_hd__dfxtp_1
X_6748__178 _6749__179/A vssd1 vssd1 vccd1 vccd1 _7622_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6690__130 _6691__131/A vssd1 vssd1 vccd1 vccd1 _7574_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput93 _5047_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[0] sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__2957_ clkbuf_0__2957_/X vssd1 vssd1 vccd1 vccd1 _6048__329/A sky130_fd_sc_hd__clkbuf_16
XFILLER_68_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4980_ _4980_/A vssd1 vssd1 vccd1 vccd1 _4980_/X sky130_fd_sc_hd__clkbuf_1
X_3931_ _3633_/X _7549_/Q _3939_/S vssd1 vssd1 vccd1 vccd1 _3932_/A sky130_fd_sc_hd__mux2_1
X_3862_ _4642_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _3878_/S sky130_fd_sc_hd__or2_4
X_6378__501 _6381__504/A vssd1 vssd1 vccd1 vccd1 _7443_/CLK sky130_fd_sc_hd__inv_2
X_5601_ _5601_/A vssd1 vssd1 vccd1 vccd1 _7084_/D sky130_fd_sc_hd__clkbuf_1
X_6581_ _6586_/B _6586_/C vssd1 vssd1 vccd1 vccd1 _6587_/B sky130_fd_sc_hd__and2_1
X_3793_ _3793_/A vssd1 vssd1 vccd1 vccd1 _7598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XCaravelHost_221 vssd1 vssd1 vccd1 vccd1 CaravelHost_221/HI partID[5] sky130_fd_sc_hd__conb_1
XCaravelHost_210 vssd1 vssd1 vccd1 vccd1 CaravelHost_210/HI manufacturerID[2] sky130_fd_sc_hd__conb_1
XCaravelHost_232 vssd1 vssd1 vccd1 vccd1 partID[2] CaravelHost_232/LO sky130_fd_sc_hd__conb_1
X_5463_ _6462_/A _5448_/X _5449_/X _5462_/X vssd1 vssd1 vccd1 vccd1 _5463_/X sky130_fd_sc_hd__a31o_1
X_7202_ _7516_/CLK _7202_/D vssd1 vssd1 vccd1 vccd1 _7202_/Q sky130_fd_sc_hd__dfxtp_2
X_4414_ _7340_/Q _4340_/X _4416_/S vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__mux2_1
X_5394_ _5385_/X _5387_/X _5393_/X _5131_/X _5161_/X vssd1 vssd1 vccd1 vccd1 _5394_/X
+ sky130_fd_sc_hd__a221o_1
X_7133_ _7133_/CLK _7133_/D vssd1 vssd1 vccd1 vccd1 _7133_/Q sky130_fd_sc_hd__dfxtp_1
X_4345_ _4345_/A vssd1 vssd1 vccd1 vccd1 _7360_/D sky130_fd_sc_hd__clkbuf_1
X_6014__301 _6017__304/A vssd1 vssd1 vccd1 vccd1 _7227_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4276_ _4276_/A vssd1 vssd1 vccd1 vccd1 _7387_/D sky130_fd_sc_hd__clkbuf_1
X_7064_ _7088_/CLK _7064_/D vssd1 vssd1 vccd1 vccd1 _7064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6970__2 _5499_/A vssd1 vssd1 vccd1 vccd1 _7712_/CLK sky130_fd_sc_hd__inv_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6623__78 _6624__79/A vssd1 vssd1 vccd1 vccd1 _7521_/CLK sky130_fd_sc_hd__inv_2
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6917_ _6917_/A _6923_/B vssd1 vssd1 vccd1 vccd1 _6918_/A sky130_fd_sc_hd__and2_1
XFILLER_50_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6848_ _6863_/D vssd1 vssd1 vccd1 vccd1 _6857_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6779_ _6779_/A _6779_/B _6779_/C _6779_/D vssd1 vssd1 vccd1 vccd1 _6878_/D sky130_fd_sc_hd__or4_4
X_6279__421 _6282__424/A vssd1 vssd1 vccd1 vccd1 _7363_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__3087_ clkbuf_0__3087_/X vssd1 vssd1 vccd1 vccd1 _6317__452/A sky130_fd_sc_hd__clkbuf_16
X_6373__497 _6373__497/A vssd1 vssd1 vccd1 vccd1 _7439_/CLK sky130_fd_sc_hd__inv_2
X_4130_ _4130_/A vssd1 vssd1 vccd1 vccd1 _7444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4061_ _4061_/A vssd1 vssd1 vccd1 vccd1 _7471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _4963_/A vssd1 vssd1 vccd1 vccd1 _4963_/X sky130_fd_sc_hd__clkbuf_1
X_6697__136 _6698__137/A vssd1 vssd1 vccd1 vccd1 _7580_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3914_ _3914_/A vssd1 vssd1 vccd1 vccd1 _3914_/X sky130_fd_sc_hd__buf_4
X_7682_ _7682_/CLK _7682_/D vssd1 vssd1 vccd1 vccd1 _7682_/Q sky130_fd_sc_hd__dfxtp_1
X_6633_ _6651_/A vssd1 vssd1 vccd1 vccd1 _6633_/X sky130_fd_sc_hd__buf_1
X_4894_ _4837_/X _7074_/Q _4898_/S vssd1 vssd1 vccd1 vccd1 _4895_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3845_ _3845_/A vssd1 vssd1 vccd1 vccd1 _7581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3776_ _4660_/A _3797_/C vssd1 vssd1 vccd1 vccd1 _3792_/S sky130_fd_sc_hd__nand2_2
X_6564_ _7505_/Q _6576_/D vssd1 vssd1 vccd1 vccd1 _6566_/B sky130_fd_sc_hd__or2_1
X_5515_ _7080_/Q _5590_/A _5515_/C vssd1 vssd1 vccd1 vccd1 _7044_/D sky130_fd_sc_hd__nor3_1
X_6495_ _6479_/X _6480_/Y _6491_/X _6505_/B _6505_/A vssd1 vssd1 vccd1 vccd1 _6495_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_118_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5446_ _5438_/X _7186_/Q _5443_/X _5445_/X vssd1 vssd1 vccd1 vccd1 _5446_/X sky130_fd_sc_hd__o22a_1
XFILLER_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5377_ _5591_/B vssd1 vssd1 vccd1 vccd1 _5494_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_113_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7116_ _7116_/CLK _7116_/D vssd1 vssd1 vccd1 vccd1 _7116_/Q sky130_fd_sc_hd__dfxtp_1
X_4328_ _7326_/Q vssd1 vssd1 vccd1 vccd1 _4328_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4259_ _4258_/X _7393_/Q _4262_/S vssd1 vssd1 vccd1 vccd1 _4260_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7047_ _7047_/CLK _7047_/D vssd1 vssd1 vccd1 vccd1 _7047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5693__249 _5693__249/A vssd1 vssd1 vccd1 vccd1 _7143_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__2959_ _6055_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2959_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2725_ clkbuf_0__2725_/X vssd1 vssd1 vccd1 vccd1 _5744__289/A sky130_fd_sc_hd__clkbuf_16
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3422_ clkbuf_0__3422_/X vssd1 vssd1 vccd1 vccd1 _6967__53/A sky130_fd_sc_hd__clkbuf_16
X_3630_ _3546_/X _7691_/Q _3630_/S vssd1 vssd1 vccd1 vccd1 _3631_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__3284_ clkbuf_0__3284_/X vssd1 vssd1 vccd1 vccd1 _6718__154/A sky130_fd_sc_hd__clkbuf_16
X_3561_ _3570_/C _4396_/A _3560_/Y vssd1 vssd1 vccd1 vccd1 _5230_/A sky130_fd_sc_hd__o21a_1
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5300_ _7133_/Q _7056_/Q _7048_/Q _7269_/Q _4374_/A _5299_/X vssd1 vssd1 vccd1 vccd1
+ _5300_/X sky130_fd_sc_hd__mux4_1
X_3492_ _4466_/C _4466_/D _4466_/B vssd1 vssd1 vccd1 vccd1 _3493_/B sky130_fd_sc_hd__mux2_1
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5231_ _5231_/A _5188_/A vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__or2b_1
XFILLER_69_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5162_ _5131_/X _5143_/X _5150_/X _5159_/X _5161_/X vssd1 vssd1 vccd1 vccd1 _5162_/X
+ sky130_fd_sc_hd__a221o_1
X_5093_ _7199_/Q _5104_/B vssd1 vssd1 vccd1 vccd1 _5094_/A sky130_fd_sc_hd__and2_1
X_4113_ _4112_/X _7450_/Q _4119_/S vssd1 vssd1 vccd1 vccd1 _4114_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4044_ _3905_/X _7478_/Q _4050_/S vssd1 vssd1 vccd1 vccd1 _4045_/A sky130_fd_sc_hd__mux2_1
X_6705__143 _6706__144/A vssd1 vssd1 vccd1 vccd1 _7587_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5995_ _5993_/X _5994_/X _5995_/S vssd1 vssd1 vccd1 vccd1 _5995_/X sky130_fd_sc_hd__mux2_2
XFILLER_52_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4946_ _3810_/X _7039_/Q _4946_/S vssd1 vssd1 vccd1 vccd1 _4947_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4877_ _4877_/A vssd1 vssd1 vccd1 vccd1 _7108_/D sky130_fd_sc_hd__clkbuf_1
X_7665_ _7727_/CLK _7665_/D vssd1 vssd1 vccd1 vccd1 _7665_/Q sky130_fd_sc_hd__dfxtp_1
X_7596_ _7596_/CLK _7596_/D vssd1 vssd1 vccd1 vccd1 _7596_/Q sky130_fd_sc_hd__dfxtp_1
X_3828_ _3735_/X _7588_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3829_/A sky130_fd_sc_hd__mux2_1
X_6616_ _6616_/A vssd1 vssd1 vccd1 vccd1 _7515_/D sky130_fd_sc_hd__clkbuf_1
X_6241__394 _6241__394/A vssd1 vssd1 vccd1 vccd1 _7334_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6547_ _7502_/Q vssd1 vssd1 vccd1 vccd1 _6553_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3759_ _3774_/S vssd1 vssd1 vccd1 vccd1 _3768_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_3_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6478_ _7504_/Q vssd1 vssd1 vccd1 vccd1 _6562_/A sky130_fd_sc_hd__clkbuf_1
X_5429_ _7161_/Q _7153_/Q _5429_/S vssd1 vssd1 vccd1 vccd1 _5429_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_1 _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3089_ _6326_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3089_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6027__311 _6027__311/A vssd1 vssd1 vccd1 vccd1 _7237_/CLK sky130_fd_sc_hd__inv_2
X_6324__458 _6325__459/A vssd1 vssd1 vccd1 vccd1 _7400_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7088_/CLK sky130_fd_sc_hd__clkbuf_8
Xclkbuf_1_1__f__2708_ clkbuf_0__2708_/X vssd1 vssd1 vccd1 vccd1 _5662__224/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4800_ _7138_/Q _4584_/A _4800_/S vssd1 vssd1 vccd1 vccd1 _4801_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5780_ _5024_/A _7200_/Q _5782_/S vssd1 vssd1 vccd1 vccd1 _5781_/A sky130_fd_sc_hd__mux2_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4731_ _4731_/A vssd1 vssd1 vccd1 vccd1 _7170_/D sky130_fd_sc_hd__clkbuf_1
X_4662_ _3794_/X _7233_/Q _4670_/S vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__mux2_1
X_7450_ _7450_/CLK _7450_/D vssd1 vssd1 vccd1 vccd1 _7450_/Q sky130_fd_sc_hd__dfxtp_1
X_6401_ _6413_/A vssd1 vssd1 vccd1 vccd1 _6401_/X sky130_fd_sc_hd__buf_1
X_3613_ _3861_/C _3796_/C _4606_/A _3822_/A vssd1 vssd1 vccd1 vccd1 _4660_/A sky130_fd_sc_hd__and4b_4
X_4593_ _4593_/A vssd1 vssd1 vccd1 vccd1 _7264_/D sky130_fd_sc_hd__clkbuf_1
X_7381_ _7381_/CLK _7381_/D vssd1 vssd1 vccd1 vccd1 _7381_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__3267_ clkbuf_0__3267_/X vssd1 vssd1 vccd1 vccd1 _6651_/A sky130_fd_sc_hd__clkbuf_16
X_3544_ _3544_/A vssd1 vssd1 vccd1 vccd1 _7708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3475_ _3822_/C vssd1 vssd1 vccd1 vccd1 _3861_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5214_ _5363_/A _5212_/X _5413_/A vssd1 vssd1 vccd1 vccd1 _5214_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5145_ _5418_/A vssd1 vssd1 vccd1 vccd1 _5289_/A sky130_fd_sc_hd__clkbuf_2
X_5076_ _5076_/A vssd1 vssd1 vccd1 vccd1 _5076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4027_ _3908_/X _7485_/Q _4031_/S vssd1 vssd1 vccd1 vccd1 _4028_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _5976_/X _5977_/X _5998_/S vssd1 vssd1 vccd1 vccd1 _5978_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ _4929_/A vssd1 vssd1 vccd1 vccd1 _7048_/D sky130_fd_sc_hd__clkbuf_1
X_7717_ _7722_/CLK _7717_/D vssd1 vssd1 vccd1 vccd1 _7717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7648_ _7655_/CLK _7648_/D vssd1 vssd1 vccd1 vccd1 _7648_/Q sky130_fd_sc_hd__dfxtp_1
X_7579_ _7579_/CLK _7579_/D vssd1 vssd1 vccd1 vccd1 _7579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6330__462 _6332__464/A vssd1 vssd1 vccd1 vccd1 _7404_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__3052_ clkbuf_0__3052_/X vssd1 vssd1 vccd1 vccd1 _6182__364/A sky130_fd_sc_hd__clkbuf_16
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5901_ _5896_/X _5899_/X _5901_/S vssd1 vssd1 vccd1 vccd1 _5902_/B sky130_fd_sc_hd__mux2_1
XFILLER_53_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6881_ _7656_/Q _6893_/B _6879_/Y _6880_/X vssd1 vssd1 vccd1 vccd1 _7656_/D sky130_fd_sc_hd__o211a_1
X_5650__214 _5650__214/A vssd1 vssd1 vccd1 vccd1 _7108_/CLK sky130_fd_sc_hd__inv_2
X_5832_ _5832_/A _5832_/B vssd1 vssd1 vccd1 vccd1 _5832_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5763_ _5763_/A vssd1 vssd1 vccd1 vccd1 _7192_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7502_ _7652_/CLK _7502_/D vssd1 vssd1 vccd1 vccd1 _7502_/Q sky130_fd_sc_hd__dfxtp_1
X_4714_ _4802_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4730_/S sky130_fd_sc_hd__or2_2
X_5694_ _5700_/A vssd1 vssd1 vccd1 vccd1 _5694_/X sky130_fd_sc_hd__buf_1
X_4645_ _4645_/A vssd1 vssd1 vccd1 vccd1 _7241_/D sky130_fd_sc_hd__clkbuf_1
X_7433_ _7433_/CLK _7433_/D vssd1 vssd1 vccd1 vccd1 _7433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4576_ _4575_/X _7269_/Q _4576_/S vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__mux2_1
X_7364_ _7364_/CLK _7364_/D vssd1 vssd1 vccd1 vccd1 _7364_/Q sky130_fd_sc_hd__dfxtp_1
X_3527_ _3526_/X _7712_/Q _3535_/S vssd1 vssd1 vccd1 vccd1 _3528_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7295_ _7295_/CLK _7295_/D vssd1 vssd1 vccd1 vccd1 _7295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6177_ _6195_/A vssd1 vssd1 vccd1 vccd1 _6177_/X sky130_fd_sc_hd__buf_1
X_5128_ _5232_/A _5380_/A _5380_/B _5380_/C vssd1 vssd1 vccd1 vccd1 _5441_/D sky130_fd_sc_hd__nor4_2
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5059_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5068_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6956__44 _6956__44/A vssd1 vssd1 vccd1 vccd1 _7700_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6174__358 _6175__359/A vssd1 vssd1 vccd1 vccd1 _7288_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4430_ _4229_/X _7333_/Q _4434_/S vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__3104_ clkbuf_0__3104_/X vssd1 vssd1 vccd1 vccd1 _6403__521/A sky130_fd_sc_hd__clkbuf_16
X_6337__468 _6337__468/A vssd1 vssd1 vccd1 vccd1 _7410_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6100_ _7650_/Q _6163_/A _6492_/C vssd1 vssd1 vccd1 vccd1 _6100_/Y sky130_fd_sc_hd__nand3b_1
X_4361_ _6272_/C _4361_/B _4361_/C vssd1 vssd1 vccd1 vccd1 _4362_/A sky130_fd_sc_hd__and3_1
X_4292_ _4292_/A vssd1 vssd1 vccd1 vccd1 _7380_/D sky130_fd_sc_hd__clkbuf_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7080_ _5496_/A _7080_/D vssd1 vssd1 vccd1 vccd1 _7080_/Q sky130_fd_sc_hd__dfxtp_1
X_6031_ _6031_/A vssd1 vssd1 vccd1 vccd1 _6031_/X sky130_fd_sc_hd__buf_1
XFILLER_100_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6864_ _6864_/A _6905_/B _6870_/C vssd1 vssd1 vccd1 vccd1 _6864_/X sky130_fd_sc_hd__or3_1
XFILLER_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5815_ _5869_/A vssd1 vssd1 vccd1 vccd1 _5855_/A sky130_fd_sc_hd__inv_2
XFILLER_50_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6795_ input1/X _6803_/B _6781_/X _6794_/X vssd1 vssd1 vccd1 vccd1 _6795_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4628_ _4243_/X _7248_/Q _4634_/S vssd1 vssd1 vccd1 vccd1 _4629_/A sky130_fd_sc_hd__mux2_1
X_7416_ _7416_/CLK _7416_/D vssd1 vssd1 vccd1 vccd1 _7416_/Q sky130_fd_sc_hd__dfxtp_1
X_4559_ _4559_/A vssd1 vssd1 vccd1 vccd1 _7277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7347_ _7347_/CLK _7347_/D vssd1 vssd1 vccd1 vccd1 _7347_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_103_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7278_ _7278_/CLK _7278_/D vssd1 vssd1 vccd1 vccd1 _7278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6229_ _7665_/Q _6231_/B vssd1 vssd1 vccd1 vccd1 _6230_/A sky130_fd_sc_hd__and2_1
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6929__22 _6930__23/A vssd1 vssd1 vccd1 vccd1 _7678_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6180__362 _6180__362/A vssd1 vssd1 vccd1 vccd1 _7292_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput94 _5069_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[10] sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__2956_ clkbuf_0__2956_/X vssd1 vssd1 vccd1 vccd1 _6041__323/A sky130_fd_sc_hd__clkbuf_16
X_5720__270 _5723__273/A vssd1 vssd1 vccd1 vccd1 _7164_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3930_ _3945_/S vssd1 vssd1 vccd1 vccd1 _3939_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6640__90 _6642__92/A vssd1 vssd1 vccd1 vccd1 _7534_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3861_ _3861_/A _6233_/A _3861_/C _3796_/C vssd1 vssd1 vccd1 vccd1 _4642_/A sky130_fd_sc_hd__or4b_4
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3792_ _3753_/X _7598_/Q _3792_/S vssd1 vssd1 vccd1 vccd1 _3793_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5600_ _7084_/Q _5057_/A _5602_/S vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6580_ _6578_/X _6579_/Y _6607_/A vssd1 vssd1 vccd1 vccd1 _7507_/D sky130_fd_sc_hd__a21oi_1
X_6950__39 _6950__39/A vssd1 vssd1 vccd1 vccd1 _7695_/CLK sky130_fd_sc_hd__inv_2
XCaravelHost_200 vssd1 vssd1 vccd1 vccd1 CaravelHost_200/HI core0Index[7] sky130_fd_sc_hd__conb_1
XCaravelHost_211 vssd1 vssd1 vccd1 vccd1 CaravelHost_211/HI manufacturerID[3] sky130_fd_sc_hd__conb_1
XCaravelHost_222 vssd1 vssd1 vccd1 vccd1 CaravelHost_222/HI partID[7] sky130_fd_sc_hd__conb_1
XCaravelHost_233 vssd1 vssd1 vccd1 vccd1 partID[4] CaravelHost_233/LO sky130_fd_sc_hd__conb_1
X_5462_ _5458_/X _7191_/Q _5450_/X input7/X vssd1 vssd1 vccd1 vccd1 _5462_/X sky130_fd_sc_hd__a22o_1
X_7201_ _7525_/CLK _7201_/D vssd1 vssd1 vccd1 vccd1 _7201_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5393_ _5264_/X _5388_/X _5390_/X _5392_/X vssd1 vssd1 vccd1 vccd1 _5393_/X sky130_fd_sc_hd__o22a_1
X_4413_ _4413_/A vssd1 vssd1 vccd1 vccd1 _7341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7132_ _7132_/CLK _7132_/D vssd1 vssd1 vccd1 vccd1 _7132_/Q sky130_fd_sc_hd__dfxtp_1
X_4344_ _7360_/Q _4343_/X _4344_/S vssd1 vssd1 vccd1 vccd1 _4345_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7063_ _7088_/CLK _7063_/D vssd1 vssd1 vccd1 vccd1 _7063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4275_ _7387_/Q _3594_/X _4275_/S vssd1 vssd1 vccd1 vccd1 _4276_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5576__207 _5576__207/A vssd1 vssd1 vccd1 vccd1 _7075_/CLK sky130_fd_sc_hd__inv_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ _6916_/A vssd1 vssd1 vccd1 vccd1 _7670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6847_ _7649_/Q _7648_/Q _6847_/C _6847_/D vssd1 vssd1 vccd1 vccd1 _6863_/D sky130_fd_sc_hd__and4_1
XFILLER_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_13_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7674_/CLK sky130_fd_sc_hd__clkbuf_8
X_6778_ _6778_/A _6778_/B _6778_/C vssd1 vssd1 vccd1 vccd1 _6779_/D sky130_fd_sc_hd__or3_1
XFILLER_23_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__3086_ clkbuf_0__3086_/X vssd1 vssd1 vccd1 vccd1 _6313__449/A sky130_fd_sc_hd__clkbuf_16
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4060_ _3899_/X _7471_/Q _4068_/S vssd1 vssd1 vccd1 vccd1 _4061_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6187__368 _6188__369/A vssd1 vssd1 vccd1 vccd1 _7298_/CLK sky130_fd_sc_hd__inv_2
X_4962_ _5642_/A _4966_/B vssd1 vssd1 vccd1 vccd1 _4963_/A sky130_fd_sc_hd__and2_1
X_6701_ _6701_/A vssd1 vssd1 vccd1 vccd1 _6701_/X sky130_fd_sc_hd__buf_1
X_3913_ _3913_/A vssd1 vssd1 vccd1 vccd1 _7554_/D sky130_fd_sc_hd__clkbuf_1
X_7681_ _7681_/CLK _7681_/D vssd1 vssd1 vccd1 vccd1 _7681_/Q sky130_fd_sc_hd__dfxtp_1
X_4893_ _4893_/A vssd1 vssd1 vccd1 vccd1 _7075_/D sky130_fd_sc_hd__clkbuf_1
X_3844_ _3730_/X _7581_/Q _3852_/S vssd1 vssd1 vccd1 vccd1 _3845_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3775_ _3775_/A vssd1 vssd1 vccd1 vccd1 _7606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6563_ _6560_/X _6562_/X _6539_/X vssd1 vssd1 vccd1 vccd1 _7504_/D sky130_fd_sc_hd__o21a_1
XFILLER_118_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5727__276 _5728__277/A vssd1 vssd1 vccd1 vccd1 _7170_/CLK sky130_fd_sc_hd__inv_2
X_5514_ _5102_/C _5513_/X _5469_/A vssd1 vssd1 vccd1 vccd1 _5515_/C sky130_fd_sc_hd__a21oi_1
X_5582__211 _5650__214/A vssd1 vssd1 vccd1 vccd1 _7079_/CLK sky130_fd_sc_hd__inv_2
X_6494_ _6163_/A _6492_/C _6586_/B vssd1 vssd1 vccd1 vccd1 _6505_/A sky130_fd_sc_hd__a21oi_1
XFILLER_105_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5445_ _5469_/A _7275_/Q _6234_/B _5381_/Y _5444_/X vssd1 vssd1 vccd1 vccd1 _5445_/X
+ sky130_fd_sc_hd__a41o_1
X_7115_ _7115_/CLK _7115_/D vssd1 vssd1 vccd1 vccd1 _7115_/Q sky130_fd_sc_hd__dfxtp_2
X_5376_ _5376_/A vssd1 vssd1 vccd1 vccd1 _5376_/X sky130_fd_sc_hd__buf_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4327_ _4327_/A vssd1 vssd1 vccd1 vccd1 _7366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4258_ _7668_/Q vssd1 vssd1 vccd1 vccd1 _4258_/X sky130_fd_sc_hd__clkbuf_2
X_7046_ _7046_/CLK _7046_/D vssd1 vssd1 vccd1 vccd1 _7046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4189_ _4115_/X _7417_/Q _4191_/S vssd1 vssd1 vccd1 vccd1 _4190_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__2958_ _6049_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2958_/X sky130_fd_sc_hd__clkbuf_16
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2724_ clkbuf_0__2724_/X vssd1 vssd1 vccd1 vccd1 _6018_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3421_ clkbuf_0__3421_/X vssd1 vssd1 vccd1 vccd1 _6962__49/A sky130_fd_sc_hd__clkbuf_16
XFILLER_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3283_ clkbuf_0__3283_/X vssd1 vssd1 vccd1 vccd1 _6710__147/A sky130_fd_sc_hd__clkbuf_16
X_3560_ _3927_/A _7348_/Q vssd1 vssd1 vccd1 vccd1 _3560_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_115_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3491_ _7316_/Q _7311_/Q vssd1 vssd1 vccd1 vccd1 _4466_/B sky130_fd_sc_hd__xnor2_1
X_5230_ _5230_/A _5230_/B _5230_/C _5230_/D vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__or4_1
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5161_ _5161_/A vssd1 vssd1 vccd1 vccd1 _5161_/X sky130_fd_sc_hd__clkbuf_2
X_5092_ _5092_/A vssd1 vssd1 vccd1 vccd1 _5104_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4112_ _7669_/Q vssd1 vssd1 vccd1 vccd1 _4112_/X sky130_fd_sc_hd__buf_2
X_4043_ _4043_/A vssd1 vssd1 vccd1 vccd1 _7479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5994_ _7589_/Q _7581_/Q _7573_/Q _7487_/Q _5912_/X _5908_/X vssd1 vssd1 vccd1 vccd1
+ _5994_/X sky130_fd_sc_hd__mux4_1
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4945_ _4945_/A vssd1 vssd1 vccd1 vccd1 _7040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4876_ _4837_/X _7108_/Q _4880_/S vssd1 vssd1 vccd1 vccd1 _4877_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7664_ _7727_/CLK _7664_/D vssd1 vssd1 vccd1 vccd1 _7664_/Q sky130_fd_sc_hd__dfxtp_1
X_3827_ _3827_/A vssd1 vssd1 vccd1 vccd1 _7589_/D sky130_fd_sc_hd__clkbuf_1
X_7595_ _7595_/CLK _7595_/D vssd1 vssd1 vccd1 vccd1 _7595_/Q sky130_fd_sc_hd__dfxtp_1
X_6615_ _6615_/A _6615_/B _6615_/C vssd1 vssd1 vccd1 vccd1 _6616_/A sky130_fd_sc_hd__and3_1
XFILLER_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6546_ _6544_/X _6545_/X _6539_/X vssd1 vssd1 vccd1 vccd1 _7501_/D sky130_fd_sc_hd__o21a_1
X_3758_ _4846_/A _4821_/A vssd1 vssd1 vccd1 vccd1 _3774_/S sky130_fd_sc_hd__or2_4
X_3689_ _3689_/A vssd1 vssd1 vccd1 vccd1 _7675_/D sky130_fd_sc_hd__clkbuf_1
X_6477_ _6483_/B _6483_/C _6483_/A vssd1 vssd1 vccd1 vccd1 _6507_/C sky130_fd_sc_hd__a21o_1
X_5428_ _4396_/A _7145_/Q _5427_/X vssd1 vssd1 vccd1 vccd1 _5428_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5359_ _7688_/Q _7611_/Q _5391_/S vssd1 vssd1 vccd1 vccd1 _5360_/B sky130_fd_sc_hd__mux2_1
XFILLER_101_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_2 _3549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7029_ _7029_/A vssd1 vssd1 vccd1 vccd1 _7730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3088_ _6320_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3088_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_55_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2707_ clkbuf_0__2707_/X vssd1 vssd1 vccd1 vccd1 _5655__218/A sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__2638_ clkbuf_0__2638_/X vssd1 vssd1 vccd1 vccd1 _5532__201/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4584_/X _7170_/Q _4730_/S vssd1 vssd1 vccd1 vccd1 _4731_/A sky130_fd_sc_hd__mux2_1
X_4661_ _4676_/S vssd1 vssd1 vccd1 vccd1 _4670_/S sky130_fd_sc_hd__buf_2
XFILLER_119_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7380_ _7380_/CLK _7380_/D vssd1 vssd1 vccd1 vccd1 _7380_/Q sky130_fd_sc_hd__dfxtp_1
X_3612_ _6915_/A _3513_/X _5535_/B vssd1 vssd1 vccd1 vccd1 _4606_/A sky130_fd_sc_hd__a21oi_4
X_4592_ _4243_/X _7264_/Q _4598_/S vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__3266_ clkbuf_0__3266_/X vssd1 vssd1 vccd1 vccd1 _6624__79/A sky130_fd_sc_hd__clkbuf_16
X_3543_ _3542_/X _7708_/Q _3547_/S vssd1 vssd1 vccd1 vccd1 _3544_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3474_ _7315_/Q vssd1 vssd1 vccd1 vccd1 _3822_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6262_ _6277_/A vssd1 vssd1 vccd1 vccd1 _6262_/X sky130_fd_sc_hd__buf_1
X_5213_ _5213_/A vssd1 vssd1 vccd1 vccd1 _5413_/A sky130_fd_sc_hd__buf_2
XFILLER_69_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5144_ _5262_/A vssd1 vssd1 vccd1 vccd1 _5418_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5075_ _5075_/A _5079_/B vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__and2_1
XFILLER_96_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4026_ _4026_/A vssd1 vssd1 vccd1 vccd1 _7486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5977_ _7248_/Q _7232_/Q _7478_/Q _7470_/Q _5860_/X _5870_/X vssd1 vssd1 vccd1 vccd1
+ _5977_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4928_ _7048_/Q _4575_/A _4928_/S vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__mux2_1
X_7716_ _7732_/CLK _7716_/D vssd1 vssd1 vccd1 vccd1 _7716_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2726_ _5745_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2726_/X sky130_fd_sc_hd__clkbuf_16
X_7647_ _7655_/CLK _7647_/D vssd1 vssd1 vccd1 vccd1 _7647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4859_/A vssd1 vssd1 vccd1 vccd1 _7116_/D sky130_fd_sc_hd__clkbuf_1
X_7578_ _7578_/CLK _7578_/D vssd1 vssd1 vccd1 vccd1 _7578_/Q sky130_fd_sc_hd__dfxtp_1
X_6529_ _6541_/C vssd1 vssd1 vccd1 vccd1 _6529_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6654__102 _6655__103/A vssd1 vssd1 vccd1 vccd1 _7546_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__3051_ clkbuf_0__3051_/X vssd1 vssd1 vccd1 vccd1 _6195_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6647__96 _6647__96/A vssd1 vssd1 vccd1 vccd1 _7540_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6266__413 _6267__414/A vssd1 vssd1 vccd1 vccd1 _7353_/CLK sky130_fd_sc_hd__inv_2
X_5900_ _5929_/A vssd1 vssd1 vccd1 vccd1 _5901_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6880_ _6886_/A vssd1 vssd1 vccd1 vccd1 _6880_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5831_ _3485_/Y _5821_/X _5825_/X _5830_/X vssd1 vssd1 vccd1 vccd1 _5832_/B sky130_fd_sc_hd__a31o_1
XFILLER_62_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5762_ _5006_/A _7192_/Q _5764_/S vssd1 vssd1 vccd1 vccd1 _5763_/A sky130_fd_sc_hd__mux2_1
X_4713_ _4713_/A vssd1 vssd1 vccd1 vccd1 _7178_/D sky130_fd_sc_hd__clkbuf_1
X_7501_ _7510_/CLK _7501_/D vssd1 vssd1 vccd1 vccd1 _7501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4644_ _4238_/X _7241_/Q _4652_/S vssd1 vssd1 vccd1 vccd1 _4645_/A sky130_fd_sc_hd__mux2_1
X_7432_ _7432_/CLK _7432_/D vssd1 vssd1 vccd1 vccd1 _7432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4575_ _4575_/A vssd1 vssd1 vccd1 vccd1 _4575_/X sky130_fd_sc_hd__clkbuf_4
X_7363_ _7363_/CLK _7363_/D vssd1 vssd1 vccd1 vccd1 _7363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3526_ _3908_/A vssd1 vssd1 vccd1 vccd1 _3526_/X sky130_fd_sc_hd__buf_2
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6314_ _6320_/A vssd1 vssd1 vccd1 vccd1 _6314_/X sky130_fd_sc_hd__buf_1
X_7294_ _7294_/CLK _7294_/D vssd1 vssd1 vccd1 vccd1 _7294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6176_ _6207_/A vssd1 vssd1 vccd1 vccd1 _6176_/X sky130_fd_sc_hd__buf_1
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5127_ _5183_/C vssd1 vssd1 vccd1 vccd1 _5380_/C sky130_fd_sc_hd__clkbuf_2
X_5058_ _5058_/A vssd1 vssd1 vccd1 vccd1 _5058_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4009_ _7493_/Q _3588_/X _4013_/S vssd1 vssd1 vccd1 vccd1 _4010_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6718__154 _6718__154/A vssd1 vssd1 vccd1 vccd1 _7598_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2709_ _5663_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2709_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5746__290 _5803__293/A vssd1 vssd1 vccd1 vccd1 _7184_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6070__346 _6071__347/A vssd1 vssd1 vccd1 vccd1 _7272_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__3103_ clkbuf_0__3103_/X vssd1 vssd1 vccd1 vccd1 _6399__518/A sky130_fd_sc_hd__clkbuf_16
X_4360_ _4363_/A _4350_/B _3927_/A vssd1 vssd1 vccd1 vccd1 _4361_/C sky130_fd_sc_hd__a21o_1
XFILLER_112_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4291_ _4249_/X _7380_/Q _4293_/S vssd1 vssd1 vccd1 vccd1 _4292_/A sky130_fd_sc_hd__mux2_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6932_ _6932_/A vssd1 vssd1 vccd1 vccd1 _6932_/X sky130_fd_sc_hd__buf_1
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6863_ _7652_/Q _7651_/Q _6863_/C _6863_/D vssd1 vssd1 vccd1 vccd1 _6870_/C sky130_fd_sc_hd__and4_1
X_5814_ _5814_/A vssd1 vssd1 vccd1 vccd1 _5814_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6794_ _6794_/A _6794_/B vssd1 vssd1 vccd1 vccd1 _6794_/X sky130_fd_sc_hd__or2_1
X_5745_ _5745_/A vssd1 vssd1 vccd1 vccd1 _5745_/X sky130_fd_sc_hd__buf_1
XFILLER_41_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5676_ _5688_/A vssd1 vssd1 vccd1 vccd1 _5676_/X sky130_fd_sc_hd__buf_1
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4627_ _4627_/A vssd1 vssd1 vccd1 vccd1 _7249_/D sky130_fd_sc_hd__clkbuf_1
X_7415_ _7415_/CLK _7415_/D vssd1 vssd1 vccd1 vccd1 _7415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4558_ _7277_/Q _3923_/A _4558_/S vssd1 vssd1 vccd1 vccd1 _4559_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7346_ _7346_/CLK _7346_/D vssd1 vssd1 vccd1 vccd1 _7346_/Q sky130_fd_sc_hd__dfxtp_1
X_7277_ _7277_/CLK _7277_/D vssd1 vssd1 vccd1 vccd1 _7277_/Q sky130_fd_sc_hd__dfxtp_1
X_4489_ _4504_/S vssd1 vssd1 vccd1 vccd1 _4498_/S sky130_fd_sc_hd__clkbuf_2
X_3509_ _7104_/Q _7103_/Q _7081_/Q vssd1 vssd1 vccd1 vccd1 _5585_/C sky130_fd_sc_hd__o21ai_1
X_6228_ _6228_/A vssd1 vssd1 vccd1 vccd1 _7326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6159_/A _6446_/B _6159_/C vssd1 vssd1 vccd1 vccd1 _6462_/B sky130_fd_sc_hd__nor3_4
XFILLER_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2955_ clkbuf_0__2955_/X vssd1 vssd1 vccd1 vccd1 _6036__319/A sky130_fd_sc_hd__clkbuf_16
XFILLER_68_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput95 _5072_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6343__473 _6344__474/A vssd1 vssd1 vccd1 vccd1 _7415_/CLK sky130_fd_sc_hd__inv_2
X_3860_ _7316_/Q vssd1 vssd1 vccd1 vccd1 _3861_/A sky130_fd_sc_hd__inv_2
XFILLER_31_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3791_ _3791_/A vssd1 vssd1 vccd1 vccd1 _7599_/D sky130_fd_sc_hd__clkbuf_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5530_ _5573_/A vssd1 vssd1 vccd1 vccd1 _5530_/X sky130_fd_sc_hd__buf_1
XFILLER_118_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XCaravelHost_212 vssd1 vssd1 vccd1 vccd1 CaravelHost_212/HI manufacturerID[4] sky130_fd_sc_hd__conb_1
X_5461_ _7719_/Q vssd1 vssd1 vccd1 vccd1 _6462_/A sky130_fd_sc_hd__buf_4
XCaravelHost_201 vssd1 vssd1 vccd1 vccd1 CaravelHost_201/HI core1Index[1] sky130_fd_sc_hd__conb_1
XFILLER_117_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XCaravelHost_223 vssd1 vssd1 vccd1 vccd1 CaravelHost_223/HI partID[9] sky130_fd_sc_hd__conb_1
XCaravelHost_234 vssd1 vssd1 vccd1 vccd1 partID[6] CaravelHost_234/LO sky130_fd_sc_hd__conb_1
X_4412_ _7341_/Q _4337_/X _4416_/S vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__mux2_1
X_7200_ _7525_/CLK _7200_/D vssd1 vssd1 vccd1 vccd1 _7200_/Q sky130_fd_sc_hd__dfxtp_4
X_5392_ _5148_/X _5391_/X _5163_/A vssd1 vssd1 vccd1 vccd1 _5392_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6667__112 _6669__114/A vssd1 vssd1 vccd1 vccd1 _7556_/CLK sky130_fd_sc_hd__inv_2
X_7131_ _7131_/CLK _7131_/D vssd1 vssd1 vccd1 vccd1 _7131_/Q sky130_fd_sc_hd__dfxtp_1
X_4343_ _7321_/Q vssd1 vssd1 vccd1 vccd1 _4343_/X sky130_fd_sc_hd__buf_4
XFILLER_113_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4274_ _4274_/A vssd1 vssd1 vccd1 vccd1 _7388_/D sky130_fd_sc_hd__clkbuf_1
X_7062_ _7088_/CLK _7062_/D vssd1 vssd1 vccd1 vccd1 _7062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6385__507 _6385__507/A vssd1 vssd1 vccd1 vccd1 _7449_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6915_ _6915_/A _6921_/B _6921_/C vssd1 vssd1 vccd1 vccd1 _6916_/A sky130_fd_sc_hd__and3_1
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6846_ _6846_/A vssd1 vssd1 vccd1 vccd1 _7648_/D sky130_fd_sc_hd__clkbuf_1
X_6777_ _6777_/A _6789_/A vssd1 vssd1 vccd1 vccd1 _6778_/C sky130_fd_sc_hd__xnor2_1
X_3989_ _3989_/A vssd1 vssd1 vccd1 vccd1 _7523_/D sky130_fd_sc_hd__clkbuf_1
X_6021__307 _6021__307/A vssd1 vssd1 vccd1 vccd1 _7233_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7329_ _7674_/CLK _7329_/D vssd1 vssd1 vccd1 vccd1 _7329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6286__427 _6287__428/A vssd1 vssd1 vccd1 vccd1 _7369_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__3085_ clkbuf_0__3085_/X vssd1 vssd1 vccd1 vccd1 _6304__441/A sky130_fd_sc_hd__clkbuf_16
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4961_ _4961_/A vssd1 vssd1 vccd1 vccd1 _4961_/X sky130_fd_sc_hd__clkbuf_1
X_3912_ _3911_/X _7554_/Q _3915_/S vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__mux2_1
X_7680_ _7680_/CLK _7680_/D vssd1 vssd1 vccd1 vccd1 _7680_/Q sky130_fd_sc_hd__dfxtp_1
X_4892_ _4834_/X _7075_/Q _4892_/S vssd1 vssd1 vccd1 vccd1 _4893_/A sky130_fd_sc_hd__mux2_1
X_3843_ _3858_/S vssd1 vssd1 vccd1 vccd1 _3852_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3774_ _3668_/X _7606_/Q _3774_/S vssd1 vssd1 vccd1 vccd1 _3775_/A sky130_fd_sc_hd__mux2_1
X_6562_ _6562_/A _6589_/B _6562_/C vssd1 vssd1 vccd1 vccd1 _6562_/X sky130_fd_sc_hd__and3_1
X_6391__511 _6392__512/A vssd1 vssd1 vccd1 vccd1 _7453_/CLK sky130_fd_sc_hd__inv_2
X_5513_ _7203_/Q _7202_/Q _7204_/Q _7205_/Q vssd1 vssd1 vccd1 vccd1 _5513_/X sky130_fd_sc_hd__and4_2
XFILLER_8_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6493_ _7508_/Q vssd1 vssd1 vccd1 vccd1 _6586_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5444_ _5458_/A vssd1 vssd1 vccd1 vccd1 _5444_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7114_ _7114_/CLK _7114_/D vssd1 vssd1 vccd1 vccd1 _7114_/Q sky130_fd_sc_hd__dfxtp_1
X_5375_ _5375_/A vssd1 vssd1 vccd1 vccd1 _5375_/X sky130_fd_sc_hd__buf_4
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4326_ _7366_/Q _4325_/X _4335_/S vssd1 vssd1 vccd1 vccd1 _4327_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4257_ _4257_/A vssd1 vssd1 vccd1 vccd1 _7394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7045_ _7045_/CLK _7045_/D vssd1 vssd1 vccd1 vccd1 _7045_/Q sky130_fd_sc_hd__dfxtp_1
X_4188_ _4188_/A vssd1 vssd1 vccd1 vccd1 _7418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__2957_ _6043_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2957_/X sky130_fd_sc_hd__clkbuf_16
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6829_ _7645_/Q _6833_/C _6829_/C vssd1 vssd1 vccd1 vccd1 _6835_/B sky130_fd_sc_hd__and3_1
XFILLER_23_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6253__404 _6253__404/A vssd1 vssd1 vccd1 vccd1 _7344_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2723_ clkbuf_0__2723_/X vssd1 vssd1 vccd1 vccd1 _6055_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3420_ clkbuf_0__3420_/X vssd1 vssd1 vccd1 vccd1 _6956__44/A sky130_fd_sc_hd__clkbuf_16
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__3282_ clkbuf_0__3282_/X vssd1 vssd1 vccd1 vccd1 _6704__142/A sky130_fd_sc_hd__clkbuf_16
X_3490_ _3822_/C _7310_/Q vssd1 vssd1 vccd1 vccd1 _4466_/D sky130_fd_sc_hd__or2b_1
XFILLER_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6193__373 _6194__374/A vssd1 vssd1 vccd1 vccd1 _7303_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5160_ _7351_/Q vssd1 vssd1 vccd1 vccd1 _5161_/A sky130_fd_sc_hd__inv_2
X_5091_ _5091_/A vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4111_ _4111_/A vssd1 vssd1 vccd1 vccd1 _7451_/D sky130_fd_sc_hd__clkbuf_1
X_4042_ _3899_/X _7479_/Q _4050_/S vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6429__61 _6429__61/A vssd1 vssd1 vccd1 vccd1 _7483_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _7541_/Q _7682_/Q _7698_/Q _7284_/Q _5907_/X _5905_/X vssd1 vssd1 vccd1 vccd1
+ _5993_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4944_ _3807_/X _7040_/Q _4946_/S vssd1 vssd1 vccd1 vccd1 _4945_/A sky130_fd_sc_hd__mux2_1
X_7732_ _7732_/CLK _7732_/D vssd1 vssd1 vccd1 vccd1 _7732_/Q sky130_fd_sc_hd__dfxtp_1
X_5733__281 _5736__284/A vssd1 vssd1 vccd1 vccd1 _7175_/CLK sky130_fd_sc_hd__inv_2
X_7663_ _7727_/CLK _7663_/D vssd1 vssd1 vccd1 vccd1 _7663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4875_ _4875_/A vssd1 vssd1 vccd1 vccd1 _7109_/D sky130_fd_sc_hd__clkbuf_1
X_3826_ _3730_/X _7589_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3827_/A sky130_fd_sc_hd__mux2_1
X_7594_ _7594_/CLK _7594_/D vssd1 vssd1 vccd1 vccd1 _7594_/Q sky130_fd_sc_hd__dfxtp_1
X_6614_ _6534_/A _6610_/Y _6515_/B vssd1 vssd1 vccd1 vccd1 _6615_/C sky130_fd_sc_hd__o21ai_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3757_ _4385_/A _4361_/B vssd1 vssd1 vccd1 vccd1 _4821_/A sky130_fd_sc_hd__or2_2
X_6545_ _7501_/Q _6556_/B _6562_/C vssd1 vssd1 vccd1 vccd1 _6545_/X sky130_fd_sc_hd__and3_1
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6712__149 _6712__149/A vssd1 vssd1 vccd1 vccd1 _7593_/CLK sky130_fd_sc_hd__inv_2
X_3688_ _3546_/X _7675_/Q _3688_/S vssd1 vssd1 vccd1 vccd1 _3689_/A sky130_fd_sc_hd__mux2_1
X_6476_ _6476_/A vssd1 vssd1 vccd1 vccd1 _6483_/A sky130_fd_sc_hd__inv_2
X_5427_ _7524_/Q _5285_/S _5252_/A vssd1 vssd1 vccd1 vccd1 _5427_/X sky130_fd_sc_hd__o21ba_1
XFILLER_114_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5740__285 _5743__288/A vssd1 vssd1 vccd1 vccd1 _7179_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5358_ _5358_/A vssd1 vssd1 vccd1 vccd1 _5358_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_3 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4309_ _4309_/A vssd1 vssd1 vccd1 vccd1 _7373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7028_ _7031_/A _7028_/B vssd1 vssd1 vccd1 vccd1 _7029_/A sky130_fd_sc_hd__or2_1
X_5289_ _5289_/A _5289_/B vssd1 vssd1 vccd1 vccd1 _5289_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_0__3087_ _6314_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3087_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6398__517 _6399__518/A vssd1 vssd1 vccd1 vccd1 _7459_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034__317 _6036__319/A vssd1 vssd1 vccd1 vccd1 _7243_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__2637_ clkbuf_0__2637_/X vssd1 vssd1 vccd1 vccd1 _5528__198/A sky130_fd_sc_hd__clkbuf_16
XFILLER_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6299__437 _6301__439/A vssd1 vssd1 vccd1 vccd1 _7379_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4660_ _4660_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _4676_/S sky130_fd_sc_hd__nand2_2
X_3611_ _3611_/A vssd1 vssd1 vccd1 vccd1 _5535_/B sky130_fd_sc_hd__clkbuf_4
X_4591_ _4591_/A vssd1 vssd1 vccd1 vccd1 _7265_/D sky130_fd_sc_hd__clkbuf_1
X_3542_ _3920_/A vssd1 vssd1 vccd1 vccd1 _3542_/X sky130_fd_sc_hd__clkbuf_2
X_3473_ _4095_/A _3900_/C _4095_/B vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__or3b_2
X_6261_ _6357_/A vssd1 vssd1 vccd1 vccd1 _6261_/X sky130_fd_sc_hd__buf_1
XFILLER_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5212_ _7155_/Q _7147_/Q _5362_/S vssd1 vssd1 vccd1 vccd1 _5212_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5143_ _5136_/X _5141_/X _5356_/A vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _5074_/A vssd1 vssd1 vccd1 vccd1 _5074_/X sky130_fd_sc_hd__clkbuf_1
X_4025_ _3905_/X _7486_/Q _4031_/S vssd1 vssd1 vccd1 vccd1 _4026_/A sky130_fd_sc_hd__mux2_1
X_6968__54 _6968__54/A vssd1 vssd1 vccd1 vccd1 _7710_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5976_ _7216_/Q _7042_/Q _7264_/Q _7256_/Q _5841_/X _5913_/X vssd1 vssd1 vccd1 vccd1
+ _5976_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4927_ _4927_/A vssd1 vssd1 vccd1 vccd1 _7049_/D sky130_fd_sc_hd__clkbuf_1
X_7715_ _7732_/CLK _7715_/D vssd1 vssd1 vccd1 vccd1 _7715_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2725_ _5739_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2725_/X sky130_fd_sc_hd__clkbuf_16
X_7646_ _7655_/CLK _7646_/D vssd1 vssd1 vccd1 vccd1 _7646_/Q sky130_fd_sc_hd__dfxtp_1
X_4858_ _4837_/X _7116_/Q _4862_/S vssd1 vssd1 vccd1 vccd1 _4859_/A sky130_fd_sc_hd__mux2_1
X_3809_ _3809_/A vssd1 vssd1 vccd1 vccd1 _7594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7577_ _7577_/CLK _7577_/D vssd1 vssd1 vccd1 vccd1 _7577_/Q sky130_fd_sc_hd__dfxtp_1
X_4789_ _4789_/A vssd1 vssd1 vccd1 vccd1 _7144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6528_ _7499_/Q vssd1 vssd1 vccd1 vccd1 _6541_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6459_ _7512_/Q _6459_/B vssd1 vssd1 vccd1 vccd1 _6509_/A sky130_fd_sc_hd__xnor2_1
XFILLER_106_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6423__56 _6424__57/A vssd1 vssd1 vccd1 vccd1 _7478_/CLK sky130_fd_sc_hd__inv_2
X_6406__524 _6406__524/A vssd1 vssd1 vccd1 vccd1 _7466_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6661__107 _6663__109/A vssd1 vssd1 vccd1 vccd1 _7551_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5830_ _5959_/S _5826_/X _5829_/X _5929_/A vssd1 vssd1 vccd1 vccd1 _5830_/X sky130_fd_sc_hd__o211a_1
XFILLER_62_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6307__444 _6307__444/A vssd1 vssd1 vccd1 vccd1 _7386_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5761_ _5761_/A vssd1 vssd1 vccd1 vccd1 _7191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7500_ _7652_/CLK _7500_/D vssd1 vssd1 vccd1 vccd1 _7500_/Q sky130_fd_sc_hd__dfxtp_1
X_4712_ _4584_/X _7178_/Q _4712_/S vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__mux2_1
X_7431_ _7431_/CLK _7431_/D vssd1 vssd1 vccd1 vccd1 _7431_/Q sky130_fd_sc_hd__dfxtp_1
X_4643_ _4658_/S vssd1 vssd1 vccd1 vccd1 _4652_/S sky130_fd_sc_hd__clkbuf_2
X_4574_ _4574_/A vssd1 vssd1 vccd1 vccd1 _7270_/D sky130_fd_sc_hd__clkbuf_1
X_7362_ _7362_/CLK _7362_/D vssd1 vssd1 vccd1 vccd1 _7362_/Q sky130_fd_sc_hd__dfxtp_1
X_3525_ _7672_/Q vssd1 vssd1 vccd1 vccd1 _3908_/A sky130_fd_sc_hd__buf_2
X_7293_ _7293_/CLK _7293_/D vssd1 vssd1 vccd1 vccd1 _7293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5126_ _7089_/Q _7090_/Q _5126_/C _5126_/D vssd1 vssd1 vccd1 vccd1 _5380_/A sky130_fd_sc_hd__or4_2
X_5057_ _5057_/A _5057_/B vssd1 vssd1 vccd1 vccd1 _5058_/A sky130_fd_sc_hd__and2_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4008_ _4008_/A vssd1 vssd1 vccd1 vccd1 _7494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5959_ _5957_/X _5958_/X _5959_/S vssd1 vssd1 vccd1 vccd1 _5959_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7629_ _7629_/CLK _7629_/D vssd1 vssd1 vccd1 vccd1 _7629_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2708_ _5657_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2708_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6725__159 _6725__159/A vssd1 vssd1 vccd1 vccd1 _7603_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6962__49 _6962__49/A vssd1 vssd1 vccd1 vccd1 _7705_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__3102_ clkbuf_0__3102_/X vssd1 vssd1 vccd1 vccd1 _6394__514/A sky130_fd_sc_hd__clkbuf_16
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4290_ _4290_/A vssd1 vssd1 vccd1 vccd1 _7381_/D sky130_fd_sc_hd__clkbuf_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6862_ _6876_/A vssd1 vssd1 vccd1 vccd1 _6905_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5813_ _5833_/A vssd1 vssd1 vccd1 vccd1 _5814_/A sky130_fd_sc_hd__buf_2
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5689__245 _5691__247/A vssd1 vssd1 vccd1 vccd1 _7139_/CLK sky130_fd_sc_hd__inv_2
X_6793_ _6789_/X _6791_/X _6792_/Y _6781_/A vssd1 vssd1 vccd1 vccd1 _6794_/B sky130_fd_sc_hd__o31ai_1
X_5675_ _5706_/A vssd1 vssd1 vccd1 vccd1 _5675_/X sky130_fd_sc_hd__buf_1
X_4626_ _4238_/X _7249_/Q _4634_/S vssd1 vssd1 vccd1 vccd1 _4627_/A sky130_fd_sc_hd__mux2_1
X_7414_ _7414_/CLK _7414_/D vssd1 vssd1 vccd1 vccd1 _7414_/Q sky130_fd_sc_hd__dfxtp_1
X_7345_ _7345_/CLK _7345_/D vssd1 vssd1 vccd1 vccd1 _7345_/Q sky130_fd_sc_hd__dfxtp_1
X_4557_ _4557_/A vssd1 vssd1 vccd1 vccd1 _7278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4488_ _4864_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4504_/S sky130_fd_sc_hd__or2_2
XFILLER_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3508_ _7085_/Q _7086_/Q _7087_/Q _7088_/Q vssd1 vssd1 vccd1 vccd1 _5585_/B sky130_fd_sc_hd__or4_2
X_7276_ _7732_/CLK _7276_/D vssd1 vssd1 vccd1 vccd1 _7276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6227_ _7664_/Q _6231_/B vssd1 vssd1 vccd1 vccd1 _6228_/A sky130_fd_sc_hd__and2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6158_/A _6158_/B _6458_/B vssd1 vssd1 vccd1 vccd1 _6771_/B sky130_fd_sc_hd__and3_1
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _7274_/Q vssd1 vssd1 vccd1 vccd1 _7010_/A sky130_fd_sc_hd__clkbuf_2
X_6089_ _7657_/Q _7656_/Q vssd1 vssd1 vccd1 vccd1 _6170_/C sky130_fd_sc_hd__and2_1
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2954_ clkbuf_0__2954_/X vssd1 vssd1 vccd1 vccd1 _6030__314/A sky130_fd_sc_hd__clkbuf_16
Xoutput96 _5074_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[12] sky130_fd_sc_hd__buf_2
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6935__27 _6937__29/A vssd1 vssd1 vccd1 vccd1 _7683_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ _3750_/X _7599_/Q _3792_/S vssd1 vssd1 vccd1 vccd1 _3791_/A sky130_fd_sc_hd__mux2_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5460_ _7720_/Q _5448_/X _5449_/X _5459_/X vssd1 vssd1 vccd1 vccd1 _5460_/X sky130_fd_sc_hd__a31o_1
XCaravelHost_202 vssd1 vssd1 vccd1 vccd1 CaravelHost_202/HI core1Index[2] sky130_fd_sc_hd__conb_1
XCaravelHost_224 vssd1 vssd1 vccd1 vccd1 CaravelHost_224/HI partID[12] sky130_fd_sc_hd__conb_1
XCaravelHost_235 vssd1 vssd1 vccd1 vccd1 partID[8] CaravelHost_235/LO sky130_fd_sc_hd__conb_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XCaravelHost_213 vssd1 vssd1 vccd1 vccd1 CaravelHost_213/HI manufacturerID[5] sky130_fd_sc_hd__conb_1
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4411_ _4411_/A vssd1 vssd1 vccd1 vccd1 _7342_/D sky130_fd_sc_hd__clkbuf_1
X_5391_ _7406_/Q _7390_/Q _5391_/S vssd1 vssd1 vccd1 vccd1 _5391_/X sky130_fd_sc_hd__mux2_1
X_7130_ _7130_/CLK _7130_/D vssd1 vssd1 vccd1 vccd1 _7130_/Q sky130_fd_sc_hd__dfxtp_1
X_4342_ _4342_/A vssd1 vssd1 vccd1 vccd1 _7361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4273_ _7388_/Q _3591_/X _4275_/S vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7061_ _7088_/CLK _7061_/D vssd1 vssd1 vccd1 vccd1 _7061_/Q sky130_fd_sc_hd__dfxtp_1
X_6012_ _6018_/A vssd1 vssd1 vccd1 vccd1 _6012_/X sky130_fd_sc_hd__buf_1
XFILLER_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
.ends

