magic
tech sky130A
magscale 1 2
timestamp 1650898099
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 170306 700544 170312 700596
rect 170364 700584 170370 700596
rect 180058 700584 180064 700596
rect 170364 700556 180064 700584
rect 170364 700544 170370 700556
rect 180058 700544 180064 700556
rect 180116 700544 180122 700596
rect 105446 700476 105452 700528
rect 105504 700516 105510 700528
rect 185578 700516 185584 700528
rect 105504 700488 185584 700516
rect 105504 700476 105510 700488
rect 185578 700476 185584 700488
rect 185636 700476 185642 700528
rect 535730 700476 535736 700528
rect 535788 700516 535794 700528
rect 543458 700516 543464 700528
rect 535788 700488 543464 700516
rect 535788 700476 535794 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 89162 700408 89168 700460
rect 89220 700448 89226 700460
rect 542998 700448 543004 700460
rect 89220 700420 543004 700448
rect 89220 700408 89226 700420
rect 542998 700408 543004 700420
rect 543056 700408 543062 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 543826 700380 543832 700392
rect 24360 700352 543832 700380
rect 24360 700340 24366 700352
rect 543826 700340 543832 700352
rect 543884 700340 543890 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 543918 700312 543924 700324
rect 8168 700284 543924 700312
rect 8168 700272 8174 700284
rect 543918 700272 543924 700284
rect 543976 700272 543982 700324
rect 348786 700068 348792 700120
rect 348844 700108 348850 700120
rect 349798 700108 349804 700120
rect 348844 700080 349804 700108
rect 348844 700068 348850 700080
rect 349798 700068 349804 700080
rect 349856 700068 349862 700120
rect 218974 699660 218980 699712
rect 219032 699700 219038 699712
rect 220078 699700 220084 699712
rect 219032 699672 220084 699700
rect 219032 699660 219038 699672
rect 220078 699660 220084 699672
rect 220136 699660 220142 699712
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 534350 696940 534356 696992
rect 534408 696980 534414 696992
rect 580166 696980 580172 696992
rect 534408 696952 580172 696980
rect 534408 696940 534414 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 193858 683176 193864 683188
rect 3476 683148 193864 683176
rect 3476 683136 3482 683148
rect 193858 683136 193864 683148
rect 193916 683136 193922 683188
rect 535546 683136 535552 683188
rect 535604 683176 535610 683188
rect 580166 683176 580172 683188
rect 535604 683148 580172 683176
rect 535604 683136 535610 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 545298 670732 545304 670744
rect 3568 670704 545304 670732
rect 3568 670692 3574 670704
rect 545298 670692 545304 670704
rect 545356 670692 545362 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 545206 656928 545212 656940
rect 3476 656900 545212 656928
rect 3476 656888 3482 656900
rect 545206 656888 545212 656900
rect 545264 656888 545270 656940
rect 554038 643084 554044 643136
rect 554096 643124 554102 643136
rect 580166 643124 580172 643136
rect 554096 643096 580172 643124
rect 554096 643084 554102 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 534166 630640 534172 630692
rect 534224 630680 534230 630692
rect 579982 630680 579988 630692
rect 534224 630652 579988 630680
rect 534224 630640 534230 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 544378 618304 544384 618316
rect 3568 618276 544384 618304
rect 3568 618264 3574 618276
rect 544378 618264 544384 618276
rect 544436 618264 544442 618316
rect 533338 616836 533344 616888
rect 533396 616876 533402 616888
rect 580166 616876 580172 616888
rect 533396 616848 580172 616876
rect 533396 616836 533402 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 546770 605860 546776 605872
rect 3568 605832 546776 605860
rect 3568 605820 3574 605832
rect 546770 605820 546776 605832
rect 546828 605820 546834 605872
rect 153194 599564 153200 599616
rect 153252 599604 153258 599616
rect 542630 599604 542636 599616
rect 153252 599576 542636 599604
rect 153252 599564 153258 599576
rect 542630 599564 542636 599576
rect 542688 599564 542694 599616
rect 532878 590656 532884 590708
rect 532936 590696 532942 590708
rect 580166 590696 580172 590708
rect 532936 590668 580172 590696
rect 532936 590656 532942 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 202874 579680 202880 579692
rect 3384 579652 202880 579680
rect 3384 579640 3390 579652
rect 202874 579640 202880 579652
rect 202932 579680 202938 579692
rect 546586 579680 546592 579692
rect 202932 579652 546592 579680
rect 202932 579640 202938 579652
rect 546586 579640 546592 579652
rect 546644 579640 546650 579692
rect 532786 576852 532792 576904
rect 532844 576892 532850 576904
rect 580166 576892 580172 576904
rect 532844 576864 580172 576892
rect 532844 576852 532850 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 177298 565876 177304 565888
rect 3292 565848 177304 565876
rect 3292 565836 3298 565848
rect 177298 565836 177304 565848
rect 177356 565836 177362 565888
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 546678 553432 546684 553444
rect 3384 553404 546684 553432
rect 3384 553392 3390 553404
rect 546678 553392 546684 553404
rect 546736 553392 546742 553444
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 208394 527184 208400 527196
rect 3016 527156 208400 527184
rect 3016 527144 3022 527156
rect 208394 527144 208400 527156
rect 208452 527184 208458 527196
rect 548150 527184 548156 527196
rect 208452 527156 548156 527184
rect 208452 527144 208458 527156
rect 548150 527144 548156 527156
rect 548208 527144 548214 527196
rect 531314 524424 531320 524476
rect 531372 524464 531378 524476
rect 580166 524464 580172 524476
rect 531372 524436 580172 524464
rect 531372 524424 531378 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 177390 514808 177396 514820
rect 3568 514780 177396 514808
rect 3568 514768 3574 514780
rect 177390 514768 177396 514780
rect 177448 514768 177454 514820
rect 299474 511912 299480 511964
rect 299532 511952 299538 511964
rect 300118 511952 300124 511964
rect 299532 511924 300124 511952
rect 299532 511912 299538 511924
rect 300118 511912 300124 511924
rect 300176 511912 300182 511964
rect 300118 510620 300124 510672
rect 300176 510660 300182 510672
rect 539870 510660 539876 510672
rect 300176 510632 539876 510660
rect 300176 510620 300182 510632
rect 539870 510620 539876 510632
rect 539928 510620 539934 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 547966 501004 547972 501016
rect 3108 500976 547972 501004
rect 3108 500964 3114 500976
rect 547966 500964 547972 500976
rect 548024 500964 548030 501016
rect 477494 497496 477500 497548
rect 477552 497536 477558 497548
rect 536834 497536 536840 497548
rect 477552 497508 536840 497536
rect 477552 497496 477558 497508
rect 536834 497496 536840 497508
rect 536892 497496 536898 497548
rect 282914 497428 282920 497480
rect 282972 497468 282978 497480
rect 539686 497468 539692 497480
rect 282972 497440 539692 497468
rect 282972 497428 282978 497440
rect 539686 497428 539692 497440
rect 539744 497428 539750 497480
rect 530118 484372 530124 484424
rect 530176 484412 530182 484424
rect 580166 484412 580172 484424
rect 530176 484384 580172 484412
rect 530176 484372 530182 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 531406 470568 531412 470620
rect 531464 470608 531470 470620
rect 579982 470608 579988 470620
rect 531464 470580 579988 470608
rect 531464 470568 531470 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 530578 456764 530584 456816
rect 530636 456804 530642 456816
rect 580166 456804 580172 456816
rect 530636 456776 580172 456804
rect 530636 456764 530642 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 527174 453296 527180 453348
rect 527232 453336 527238 453348
rect 535638 453336 535644 453348
rect 527232 453308 535644 453336
rect 527232 453296 527238 453308
rect 535638 453296 535644 453308
rect 535696 453296 535702 453348
rect 529658 430584 529664 430636
rect 529716 430624 529722 430636
rect 580166 430624 580172 430636
rect 529716 430596 580172 430624
rect 529716 430584 529722 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 539778 428856 539784 428868
rect 538968 428828 539784 428856
rect 412634 428748 412640 428800
rect 412692 428788 412698 428800
rect 538490 428788 538496 428800
rect 412692 428760 538496 428788
rect 412692 428748 412698 428760
rect 538490 428748 538496 428760
rect 538548 428748 538554 428800
rect 349798 428680 349804 428732
rect 349856 428720 349862 428732
rect 538968 428720 538996 428828
rect 539778 428816 539784 428828
rect 539836 428816 539842 428868
rect 541526 428788 541532 428800
rect 349856 428692 538996 428720
rect 539612 428760 541532 428788
rect 349856 428680 349862 428692
rect 220078 428612 220084 428664
rect 220136 428652 220142 428664
rect 539612 428652 539640 428760
rect 541526 428748 541532 428760
rect 541584 428748 541590 428800
rect 220136 428624 539640 428652
rect 220136 428612 220142 428624
rect 539686 428612 539692 428664
rect 539744 428652 539750 428664
rect 540514 428652 540520 428664
rect 539744 428624 540520 428652
rect 539744 428612 539750 428624
rect 540514 428612 540520 428624
rect 540572 428612 540578 428664
rect 177390 428544 177396 428596
rect 177448 428584 177454 428596
rect 548886 428584 548892 428596
rect 177448 428556 548892 428584
rect 177448 428544 177454 428556
rect 548886 428544 548892 428556
rect 548944 428544 548950 428596
rect 177298 428476 177304 428528
rect 177356 428516 177362 428528
rect 548058 428516 548064 428528
rect 177356 428488 548064 428516
rect 177356 428476 177362 428488
rect 548058 428476 548064 428488
rect 548116 428476 548122 428528
rect 3602 428408 3608 428460
rect 3660 428448 3666 428460
rect 549990 428448 549996 428460
rect 3660 428420 549996 428448
rect 3660 428408 3666 428420
rect 549990 428408 549996 428420
rect 550048 428408 550054 428460
rect 534350 427456 534356 427508
rect 534408 427496 534414 427508
rect 554038 427496 554044 427508
rect 534408 427468 554044 427496
rect 534408 427456 534414 427468
rect 554038 427456 554044 427468
rect 554096 427456 554102 427508
rect 531866 427388 531872 427440
rect 531924 427428 531930 427440
rect 580442 427428 580448 427440
rect 531924 427400 580448 427428
rect 531924 427388 531930 427400
rect 580442 427388 580448 427400
rect 580500 427388 580506 427440
rect 462314 427320 462320 427372
rect 462372 427360 462378 427372
rect 537018 427360 537024 427372
rect 462372 427332 537024 427360
rect 462372 427320 462378 427332
rect 537018 427320 537024 427332
rect 537076 427320 537082 427372
rect 397454 427252 397460 427304
rect 397512 427292 397518 427304
rect 538214 427292 538220 427304
rect 397512 427264 538220 427292
rect 397512 427252 397518 427264
rect 538214 427252 538220 427264
rect 538272 427252 538278 427304
rect 201494 427184 201500 427236
rect 201552 427224 201558 427236
rect 541158 427224 541164 427236
rect 201552 427196 541164 427224
rect 201552 427184 201558 427196
rect 541158 427184 541164 427196
rect 541216 427184 541222 427236
rect 71774 427116 71780 427168
rect 71832 427156 71838 427168
rect 543274 427156 543280 427168
rect 71832 427128 543280 427156
rect 71832 427116 71838 427128
rect 543274 427116 543280 427128
rect 543332 427116 543338 427168
rect 3694 427048 3700 427100
rect 3752 427088 3758 427100
rect 549622 427088 549628 427100
rect 3752 427060 549628 427088
rect 3752 427048 3758 427060
rect 549622 427048 549628 427060
rect 549680 427048 549686 427100
rect 364334 426368 364340 426420
rect 364392 426408 364398 426420
rect 364978 426408 364984 426420
rect 364392 426380 364984 426408
rect 364392 426368 364398 426380
rect 364978 426368 364984 426380
rect 365036 426368 365042 426420
rect 535178 425892 535184 425944
rect 535236 425932 535242 425944
rect 580258 425932 580264 425944
rect 535236 425904 580264 425932
rect 535236 425892 535242 425904
rect 580258 425892 580264 425904
rect 580316 425892 580322 425944
rect 331214 425824 331220 425876
rect 331272 425864 331278 425876
rect 539134 425864 539140 425876
rect 331272 425836 539140 425864
rect 331272 425824 331278 425836
rect 539134 425824 539140 425836
rect 539192 425824 539198 425876
rect 3510 425756 3516 425808
rect 3568 425796 3574 425808
rect 212534 425796 212540 425808
rect 3568 425768 212540 425796
rect 3568 425756 3574 425768
rect 212534 425756 212540 425768
rect 212592 425756 212598 425808
rect 266354 425756 266360 425808
rect 266412 425796 266418 425808
rect 540146 425796 540152 425808
rect 266412 425768 540152 425796
rect 266412 425756 266418 425768
rect 540146 425756 540152 425768
rect 540204 425756 540210 425808
rect 136634 425688 136640 425740
rect 136692 425728 136698 425740
rect 542354 425728 542360 425740
rect 136692 425700 542360 425728
rect 136692 425688 136698 425700
rect 542354 425688 542360 425700
rect 542412 425688 542418 425740
rect 184934 425552 184940 425604
rect 184992 425592 184998 425604
rect 185578 425592 185584 425604
rect 184992 425564 185584 425592
rect 184992 425552 184998 425564
rect 185578 425552 185584 425564
rect 185636 425552 185642 425604
rect 364978 425212 364984 425264
rect 365036 425252 365042 425264
rect 538858 425252 538864 425264
rect 365036 425224 538864 425252
rect 365036 425212 365042 425224
rect 538858 425212 538864 425224
rect 538916 425212 538922 425264
rect 212534 425144 212540 425196
rect 212592 425184 212598 425196
rect 549346 425184 549352 425196
rect 212592 425156 549352 425184
rect 212592 425144 212598 425156
rect 549346 425144 549352 425156
rect 549404 425144 549410 425196
rect 185578 425076 185584 425128
rect 185636 425116 185642 425128
rect 543090 425116 543096 425128
rect 185636 425088 543096 425116
rect 185636 425076 185642 425088
rect 543090 425076 543096 425088
rect 543148 425076 543154 425128
rect 234614 425008 234620 425060
rect 234672 425048 234678 425060
rect 235258 425048 235264 425060
rect 234672 425020 235264 425048
rect 234672 425008 234678 425020
rect 235258 425008 235264 425020
rect 235316 425008 235322 425060
rect 542998 425008 543004 425060
rect 543056 425048 543062 425060
rect 543734 425048 543740 425060
rect 543056 425020 543740 425048
rect 543056 425008 543062 425020
rect 543734 425008 543740 425020
rect 543792 425008 543798 425060
rect 532786 424668 532792 424720
rect 532844 424708 532850 424720
rect 533154 424708 533160 424720
rect 532844 424680 533160 424708
rect 532844 424668 532850 424680
rect 533154 424668 533160 424680
rect 533212 424668 533218 424720
rect 494054 424640 494060 424652
rect 489886 424612 494060 424640
rect 445018 424396 445024 424448
rect 445076 424436 445082 424448
rect 489886 424436 489914 424612
rect 494054 424600 494060 424612
rect 494112 424640 494118 424652
rect 536834 424640 536840 424652
rect 494112 424612 536840 424640
rect 494112 424600 494118 424612
rect 536834 424600 536840 424612
rect 536892 424600 536898 424652
rect 536742 424532 536748 424584
rect 536800 424572 536806 424584
rect 558914 424572 558920 424584
rect 536800 424544 558920 424572
rect 536800 424532 536806 424544
rect 558914 424532 558920 424544
rect 558972 424532 558978 424584
rect 532786 424464 532792 424516
rect 532844 424504 532850 424516
rect 580350 424504 580356 424516
rect 532844 424476 580356 424504
rect 532844 424464 532850 424476
rect 580350 424464 580356 424476
rect 580408 424464 580414 424516
rect 445076 424408 489914 424436
rect 445076 424396 445082 424408
rect 531682 424396 531688 424448
rect 531740 424436 531746 424448
rect 580534 424436 580540 424448
rect 531740 424408 580540 424436
rect 531740 424396 531746 424408
rect 580534 424396 580540 424408
rect 580592 424396 580598 424448
rect 3418 424328 3424 424380
rect 3476 424368 3482 424380
rect 198734 424368 198740 424380
rect 3476 424340 198740 424368
rect 3476 424328 3482 424340
rect 198734 424328 198740 424340
rect 198792 424328 198798 424380
rect 429194 424328 429200 424380
rect 429252 424368 429258 424380
rect 529198 424368 529204 424380
rect 429252 424340 529204 424368
rect 429252 424328 429258 424340
rect 529198 424328 529204 424340
rect 529256 424328 529262 424380
rect 235258 423920 235264 423972
rect 235316 423960 235322 423972
rect 540974 423960 540980 423972
rect 235316 423932 540980 423960
rect 235316 423920 235322 423932
rect 540974 423920 540980 423932
rect 541032 423920 541038 423972
rect 543660 423932 543872 423960
rect 198734 423852 198740 423904
rect 198792 423892 198798 423904
rect 543660 423892 543688 423932
rect 198792 423864 543688 423892
rect 543844 423892 543872 423932
rect 544378 423920 544384 423972
rect 544436 423960 544442 423972
rect 546954 423960 546960 423972
rect 544436 423932 546960 423960
rect 544436 423920 544442 423932
rect 546954 423920 546960 423932
rect 547012 423920 547018 423972
rect 546126 423892 546132 423904
rect 543844 423864 546132 423892
rect 198792 423852 198798 423864
rect 546126 423852 546132 423864
rect 546184 423852 546190 423904
rect 546678 423852 546684 423904
rect 546736 423892 546742 423904
rect 547506 423892 547512 423904
rect 546736 423864 547512 423892
rect 546736 423852 546742 423864
rect 547506 423852 547512 423864
rect 547564 423852 547570 423904
rect 179414 423784 179420 423836
rect 179472 423824 179478 423836
rect 180058 423824 180064 423836
rect 179472 423796 180064 423824
rect 179472 423784 179478 423796
rect 180058 423784 180064 423796
rect 180116 423824 180122 423836
rect 541894 423824 541900 423836
rect 180116 423796 541900 423824
rect 180116 423784 180122 423796
rect 541894 423784 541900 423796
rect 541952 423784 541958 423836
rect 543826 423784 543832 423836
rect 543884 423824 543890 423836
rect 544746 423824 544752 423836
rect 543884 423796 544752 423824
rect 543884 423784 543890 423796
rect 544746 423784 544752 423796
rect 544804 423784 544810 423836
rect 546586 423784 546592 423836
rect 546644 423824 546650 423836
rect 547138 423824 547144 423836
rect 546644 423796 547144 423824
rect 546644 423784 546650 423796
rect 547138 423784 547144 423796
rect 547196 423784 547202 423836
rect 547966 423784 547972 423836
rect 548024 423824 548030 423836
rect 548610 423824 548616 423836
rect 548024 423796 548616 423824
rect 548024 423784 548030 423796
rect 548610 423784 548616 423796
rect 548668 423784 548674 423836
rect 77938 423716 77944 423768
rect 77996 423756 78002 423768
rect 556982 423756 556988 423768
rect 77996 423728 556988 423756
rect 77996 423716 78002 423728
rect 556982 423716 556988 423728
rect 557040 423716 557046 423768
rect 4890 423648 4896 423700
rect 4948 423688 4954 423700
rect 4948 423660 540974 423688
rect 4948 423648 4954 423660
rect 530118 423580 530124 423632
rect 530176 423620 530182 423632
rect 530854 423620 530860 423632
rect 530176 423592 530860 423620
rect 530176 423580 530182 423592
rect 530854 423580 530860 423592
rect 530912 423580 530918 423632
rect 531314 423580 531320 423632
rect 531372 423620 531378 423632
rect 532050 423620 532056 423632
rect 531372 423592 532056 423620
rect 531372 423580 531378 423592
rect 532050 423580 532056 423592
rect 532108 423580 532114 423632
rect 540946 423552 540974 423660
rect 550358 423552 550364 423564
rect 540946 423524 550364 423552
rect 550358 423512 550364 423524
rect 550416 423512 550422 423564
rect 445294 423240 445300 423292
rect 445352 423280 445358 423292
rect 533522 423280 533528 423292
rect 445352 423252 533528 423280
rect 445352 423240 445358 423252
rect 533522 423240 533528 423252
rect 533580 423240 533586 423292
rect 445110 423172 445116 423224
rect 445168 423212 445174 423224
rect 535730 423212 535736 423224
rect 445168 423184 535736 423212
rect 445168 423172 445174 423184
rect 535730 423172 535736 423184
rect 535788 423212 535794 423224
rect 536742 423212 536748 423224
rect 535788 423184 536748 423212
rect 535788 423172 535794 423184
rect 536742 423172 536748 423184
rect 536800 423172 536806 423224
rect 524138 423104 524144 423156
rect 524196 423144 524202 423156
rect 547782 423144 547788 423156
rect 524196 423116 547788 423144
rect 524196 423104 524202 423116
rect 547782 423104 547788 423116
rect 547840 423104 547846 423156
rect 175918 423036 175924 423088
rect 175976 423076 175982 423088
rect 553578 423076 553584 423088
rect 175976 423048 553584 423076
rect 175976 423036 175982 423048
rect 553578 423036 553584 423048
rect 553636 423036 553642 423088
rect 4062 422968 4068 423020
rect 4120 423008 4126 423020
rect 4890 423008 4896 423020
rect 4120 422980 4896 423008
rect 4120 422968 4126 422980
rect 4890 422968 4896 422980
rect 4948 422968 4954 423020
rect 87598 422968 87604 423020
rect 87656 423008 87662 423020
rect 552198 423008 552204 423020
rect 87656 422980 552204 423008
rect 87656 422968 87662 422980
rect 552198 422968 552204 422980
rect 552256 422968 552262 423020
rect 43438 422900 43444 422952
rect 43496 422940 43502 422952
rect 551002 422940 551008 422952
rect 43496 422912 551008 422940
rect 43496 422900 43502 422912
rect 551002 422900 551008 422912
rect 551060 422900 551066 422952
rect 522942 422832 522948 422884
rect 523000 422872 523006 422884
rect 549254 422872 549260 422884
rect 523000 422844 549260 422872
rect 523000 422832 523006 422844
rect 549254 422832 549260 422844
rect 549312 422832 549318 422884
rect 522022 422764 522028 422816
rect 522080 422804 522086 422816
rect 561030 422804 561036 422816
rect 522080 422776 561036 422804
rect 522080 422764 522086 422776
rect 561030 422764 561036 422776
rect 561088 422764 561094 422816
rect 529014 422696 529020 422748
rect 529072 422736 529078 422748
rect 548518 422736 548524 422748
rect 529072 422708 548524 422736
rect 529072 422696 529078 422708
rect 548518 422696 548524 422708
rect 548576 422696 548582 422748
rect 445202 422628 445208 422680
rect 445260 422668 445266 422680
rect 534718 422668 534724 422680
rect 445260 422640 534724 422668
rect 445260 422628 445266 422640
rect 534718 422628 534724 422640
rect 534776 422668 534782 422680
rect 535178 422668 535184 422680
rect 534776 422640 535184 422668
rect 534776 422628 534782 422640
rect 535178 422628 535184 422640
rect 535236 422628 535242 422680
rect 535270 422628 535276 422680
rect 535328 422668 535334 422680
rect 558362 422668 558368 422680
rect 535328 422640 558368 422668
rect 535328 422628 535334 422640
rect 558362 422628 558368 422640
rect 558420 422628 558426 422680
rect 530486 422560 530492 422612
rect 530544 422600 530550 422612
rect 561674 422600 561680 422612
rect 530544 422572 561680 422600
rect 530544 422560 530550 422572
rect 561674 422560 561680 422572
rect 561732 422560 561738 422612
rect 352558 422492 352564 422544
rect 352616 422532 352622 422544
rect 554222 422532 554228 422544
rect 352616 422504 554228 422532
rect 352616 422492 352622 422504
rect 554222 422492 554228 422504
rect 554280 422492 554286 422544
rect 525702 422424 525708 422476
rect 525760 422464 525766 422476
rect 535362 422464 535368 422476
rect 525760 422436 535368 422464
rect 525760 422424 525766 422436
rect 535362 422424 535368 422436
rect 535420 422424 535426 422476
rect 526254 422356 526260 422408
rect 526312 422396 526318 422408
rect 538766 422396 538772 422408
rect 526312 422368 538772 422396
rect 526312 422356 526318 422368
rect 538766 422356 538772 422368
rect 538824 422356 538830 422408
rect 523770 422288 523776 422340
rect 523828 422328 523834 422340
rect 529934 422328 529940 422340
rect 523828 422300 529940 422328
rect 523828 422288 523834 422300
rect 529934 422288 529940 422300
rect 529992 422288 529998 422340
rect 550634 422288 550640 422340
rect 550692 422328 550698 422340
rect 558086 422328 558092 422340
rect 550692 422300 558092 422328
rect 550692 422288 550698 422300
rect 558086 422288 558092 422300
rect 558144 422288 558150 422340
rect 126974 421948 126980 422000
rect 127032 421988 127038 422000
rect 530762 421988 530768 422000
rect 127032 421960 530768 421988
rect 127032 421948 127038 421960
rect 530762 421948 530768 421960
rect 530820 421948 530826 422000
rect 284938 421880 284944 421932
rect 284996 421920 285002 421932
rect 529290 421920 529296 421932
rect 284996 421892 529296 421920
rect 284996 421880 285002 421892
rect 529290 421880 529296 421892
rect 529348 421880 529354 421932
rect 548518 421880 548524 421932
rect 548576 421920 548582 421932
rect 580810 421920 580816 421932
rect 548576 421892 580816 421920
rect 548576 421880 548582 421892
rect 580810 421880 580816 421892
rect 580868 421880 580874 421932
rect 527634 421812 527640 421864
rect 527692 421852 527698 421864
rect 560662 421852 560668 421864
rect 527692 421824 560668 421852
rect 527692 421812 527698 421824
rect 560662 421812 560668 421824
rect 560720 421812 560726 421864
rect 528462 421744 528468 421796
rect 528520 421784 528526 421796
rect 560754 421784 560760 421796
rect 528520 421756 560760 421784
rect 528520 421744 528526 421756
rect 560754 421744 560760 421756
rect 560812 421744 560818 421796
rect 136634 421676 136640 421728
rect 136692 421716 136698 421728
rect 532786 421716 532792 421728
rect 136692 421688 532792 421716
rect 136692 421676 136698 421688
rect 532786 421676 532792 421688
rect 532844 421676 532850 421728
rect 535362 421676 535368 421728
rect 535420 421716 535426 421728
rect 580718 421716 580724 421728
rect 535420 421688 580724 421716
rect 535420 421676 535426 421688
rect 580718 421676 580724 421688
rect 580776 421676 580782 421728
rect 3694 421608 3700 421660
rect 3752 421648 3758 421660
rect 527082 421648 527088 421660
rect 3752 421620 527088 421648
rect 3752 421608 3758 421620
rect 527082 421608 527088 421620
rect 527140 421608 527146 421660
rect 529934 421608 529940 421660
rect 529992 421648 529998 421660
rect 580534 421648 580540 421660
rect 529992 421620 580540 421648
rect 529992 421608 529998 421620
rect 580534 421608 580540 421620
rect 580592 421608 580598 421660
rect 3878 421540 3884 421592
rect 3936 421580 3942 421592
rect 550634 421580 550640 421592
rect 3936 421552 550640 421580
rect 3936 421540 3942 421552
rect 550634 421540 550640 421552
rect 550692 421540 550698 421592
rect 528922 421472 528928 421524
rect 528980 421512 528986 421524
rect 563882 421512 563888 421524
rect 528980 421484 563888 421512
rect 528980 421472 528986 421484
rect 563882 421472 563888 421484
rect 563940 421472 563946 421524
rect 528002 421404 528008 421456
rect 528060 421444 528066 421456
rect 563790 421444 563796 421456
rect 528060 421416 563796 421444
rect 528060 421404 528066 421416
rect 563790 421404 563796 421416
rect 563848 421404 563854 421456
rect 526898 421336 526904 421388
rect 526956 421376 526962 421388
rect 562410 421376 562416 421388
rect 526956 421348 562416 421376
rect 526956 421336 526962 421348
rect 562410 421336 562416 421348
rect 562468 421336 562474 421388
rect 521010 421268 521016 421320
rect 521068 421308 521074 421320
rect 560938 421308 560944 421320
rect 521068 421280 560944 421308
rect 521068 421268 521074 421280
rect 560938 421268 560944 421280
rect 560996 421268 561002 421320
rect 521562 421200 521568 421252
rect 521620 421240 521626 421252
rect 561122 421240 561128 421252
rect 521620 421212 561128 421240
rect 521620 421200 521626 421212
rect 561122 421200 561128 421212
rect 561180 421200 561186 421252
rect 520642 421132 520648 421184
rect 520700 421172 520706 421184
rect 580258 421172 580264 421184
rect 520700 421144 580264 421172
rect 520700 421132 520706 421144
rect 580258 421132 580264 421144
rect 580316 421132 580322 421184
rect 522758 421064 522764 421116
rect 522816 421104 522822 421116
rect 561214 421104 561220 421116
rect 522816 421076 561220 421104
rect 522816 421064 522822 421076
rect 561214 421064 561220 421076
rect 561272 421064 561278 421116
rect 524874 420996 524880 421048
rect 524932 421036 524938 421048
rect 562318 421036 562324 421048
rect 524932 421008 562324 421036
rect 524932 420996 524938 421008
rect 562318 420996 562324 421008
rect 562376 420996 562382 421048
rect 525242 420928 525248 420980
rect 525300 420968 525306 420980
rect 569218 420968 569224 420980
rect 525300 420940 569224 420968
rect 525300 420928 525306 420940
rect 569218 420928 569224 420940
rect 569276 420928 569282 420980
rect 529198 420860 529204 420912
rect 529256 420900 529262 420912
rect 537662 420900 537668 420912
rect 529256 420872 537668 420900
rect 529256 420860 529262 420872
rect 537662 420860 537668 420872
rect 537720 420860 537726 420912
rect 538766 420588 538772 420640
rect 538824 420628 538830 420640
rect 542722 420628 542728 420640
rect 538824 420600 542728 420628
rect 538824 420588 538830 420600
rect 542722 420588 542728 420600
rect 542780 420588 542786 420640
rect 525886 420452 525892 420504
rect 525944 420492 525950 420504
rect 539410 420492 539416 420504
rect 525944 420464 539416 420492
rect 525944 420452 525950 420464
rect 539410 420452 539416 420464
rect 539468 420452 539474 420504
rect 524506 420384 524512 420436
rect 524564 420424 524570 420436
rect 541342 420424 541348 420436
rect 524564 420396 541348 420424
rect 524564 420384 524570 420396
rect 541342 420384 541348 420396
rect 541400 420384 541406 420436
rect 541618 420384 541624 420436
rect 541676 420424 541682 420436
rect 547966 420424 547972 420436
rect 541676 420396 547972 420424
rect 541676 420384 541682 420396
rect 547966 420384 547972 420396
rect 548024 420384 548030 420436
rect 549254 420384 549260 420436
rect 549312 420424 549318 420436
rect 580350 420424 580356 420436
rect 549312 420396 580356 420424
rect 549312 420384 549318 420396
rect 580350 420384 580356 420396
rect 580408 420384 580414 420436
rect 530118 420316 530124 420368
rect 530176 420356 530182 420368
rect 546678 420356 546684 420368
rect 530176 420328 546684 420356
rect 530176 420316 530182 420328
rect 546678 420316 546684 420328
rect 546736 420316 546742 420368
rect 547782 420316 547788 420368
rect 547840 420356 547846 420368
rect 580442 420356 580448 420368
rect 547840 420328 580448 420356
rect 547840 420316 547846 420328
rect 580442 420316 580448 420328
rect 580500 420316 580506 420368
rect 530026 420248 530032 420300
rect 530084 420288 530090 420300
rect 541618 420288 541624 420300
rect 530084 420260 541624 420288
rect 530084 420248 530090 420260
rect 541618 420248 541624 420260
rect 541676 420248 541682 420300
rect 542722 420248 542728 420300
rect 542780 420288 542786 420300
rect 580626 420288 580632 420300
rect 542780 420260 580632 420288
rect 542780 420248 542786 420260
rect 580626 420248 580632 420260
rect 580684 420248 580690 420300
rect 232498 420180 232504 420232
rect 232556 420220 232562 420232
rect 553670 420220 553676 420232
rect 232556 420192 553676 420220
rect 232556 420180 232562 420192
rect 553670 420180 553676 420192
rect 553728 420180 553734 420232
rect 132494 420112 132500 420164
rect 132552 420152 132558 420164
rect 531682 420152 531688 420164
rect 132552 420124 531688 420152
rect 132552 420112 132558 420124
rect 531682 420112 531688 420124
rect 531740 420112 531746 420164
rect 539410 420112 539416 420164
rect 539468 420152 539474 420164
rect 546586 420152 546592 420164
rect 539468 420124 546592 420152
rect 539468 420112 539474 420124
rect 546586 420112 546592 420124
rect 546644 420112 546650 420164
rect 160094 420044 160100 420096
rect 160152 420084 160158 420096
rect 429194 420084 429200 420096
rect 160152 420056 429200 420084
rect 160152 420044 160158 420056
rect 429194 420044 429200 420056
rect 429252 420044 429258 420096
rect 529474 420044 529480 420096
rect 529532 420084 529538 420096
rect 562502 420084 562508 420096
rect 529532 420056 562508 420084
rect 529532 420044 529538 420056
rect 562502 420044 562508 420056
rect 562560 420044 562566 420096
rect 527358 419976 527364 420028
rect 527416 420016 527422 420028
rect 527416 419988 532694 420016
rect 527416 419976 527422 419988
rect 530026 419948 530032 419960
rect 509206 419920 530032 419948
rect 445478 419840 445484 419892
rect 445536 419880 445542 419892
rect 509206 419880 509234 419920
rect 530026 419908 530032 419920
rect 530084 419908 530090 419960
rect 532666 419948 532694 419988
rect 541342 419976 541348 420028
rect 541400 420016 541406 420028
rect 560386 420016 560392 420028
rect 541400 419988 550634 420016
rect 541400 419976 541406 419988
rect 550606 419948 550634 419988
rect 554516 419988 560392 420016
rect 554516 419948 554544 419988
rect 560386 419976 560392 419988
rect 560444 419976 560450 420028
rect 555694 419948 555700 419960
rect 532666 419920 546494 419948
rect 550606 419920 554544 419948
rect 554608 419920 555700 419948
rect 530118 419880 530124 419892
rect 445536 419852 509234 419880
rect 528296 419852 530124 419880
rect 445536 419840 445542 419852
rect 445662 419772 445668 419824
rect 445720 419812 445726 419824
rect 525886 419812 525892 419824
rect 445720 419784 525892 419812
rect 445720 419772 445726 419784
rect 525886 419772 525892 419784
rect 525944 419772 525950 419824
rect 236638 419704 236644 419756
rect 236696 419744 236702 419756
rect 528296 419744 528324 419852
rect 530118 419840 530124 419852
rect 530176 419840 530182 419892
rect 540946 419852 545896 419880
rect 528370 419772 528376 419824
rect 528428 419772 528434 419824
rect 236696 419716 528324 419744
rect 236696 419704 236702 419716
rect 193858 419636 193864 419688
rect 193916 419676 193922 419688
rect 193916 419648 509234 419676
rect 193916 419636 193922 419648
rect 509206 419608 509234 419648
rect 519814 419608 519820 419620
rect 509206 419580 519820 419608
rect 519814 419568 519820 419580
rect 519872 419568 519878 419620
rect 193214 419500 193220 419552
rect 193272 419540 193278 419552
rect 193858 419540 193864 419552
rect 193272 419512 193864 419540
rect 193272 419500 193278 419512
rect 193858 419500 193864 419512
rect 193916 419500 193922 419552
rect 514662 419500 514668 419552
rect 514720 419540 514726 419552
rect 517514 419540 517520 419552
rect 514720 419512 517520 419540
rect 514720 419500 514726 419512
rect 517514 419500 517520 419512
rect 517572 419500 517578 419552
rect 528388 419472 528416 419772
rect 528388 419444 532694 419472
rect 532666 419268 532694 419444
rect 532666 419240 536834 419268
rect 536806 419132 536834 419240
rect 540946 419132 540974 419852
rect 545206 419772 545212 419824
rect 545264 419772 545270 419824
rect 536806 419104 540974 419132
rect 519814 418956 519820 419008
rect 519872 418996 519878 419008
rect 519872 418968 524414 418996
rect 519872 418956 519878 418968
rect 524386 418928 524414 418968
rect 545224 418928 545252 419772
rect 545868 419540 545896 419852
rect 546466 419608 546494 419920
rect 547966 419840 547972 419892
rect 548024 419880 548030 419892
rect 554608 419880 554636 419920
rect 555694 419908 555700 419920
rect 555752 419908 555758 419960
rect 548024 419852 554636 419880
rect 548024 419840 548030 419852
rect 546586 419772 546592 419824
rect 546644 419772 546650 419824
rect 546678 419772 546684 419824
rect 546736 419812 546742 419824
rect 546736 419784 546816 419812
rect 546736 419772 546742 419784
rect 546604 419676 546632 419772
rect 546788 419744 546816 419784
rect 554590 419772 554596 419824
rect 554648 419772 554654 419824
rect 556706 419772 556712 419824
rect 556764 419772 556770 419824
rect 559282 419772 559288 419824
rect 559340 419812 559346 419824
rect 559926 419812 559932 419824
rect 559340 419784 559932 419812
rect 559340 419772 559346 419784
rect 559926 419772 559932 419784
rect 559984 419772 559990 419824
rect 560018 419772 560024 419824
rect 560076 419812 560082 419824
rect 560202 419812 560208 419824
rect 560076 419784 560208 419812
rect 560076 419772 560082 419784
rect 560202 419772 560208 419784
rect 560260 419772 560266 419824
rect 554608 419744 554636 419772
rect 546788 419716 554636 419744
rect 556724 419676 556752 419772
rect 546604 419648 556752 419676
rect 563698 419608 563704 419620
rect 546466 419580 563704 419608
rect 563698 419568 563704 419580
rect 563756 419568 563762 419620
rect 566458 419540 566464 419552
rect 545868 419512 566464 419540
rect 566458 419500 566464 419512
rect 566516 419500 566522 419552
rect 561674 419432 561680 419484
rect 561732 419472 561738 419484
rect 580166 419472 580172 419484
rect 561732 419444 580172 419472
rect 561732 419432 561738 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 524386 418900 545252 418928
rect 447594 416848 447600 416900
rect 447652 416888 447658 416900
rect 517514 416888 517520 416900
rect 447652 416860 517520 416888
rect 447652 416848 447658 416860
rect 517514 416848 517520 416860
rect 517572 416848 517578 416900
rect 447870 416780 447876 416832
rect 447928 416820 447934 416832
rect 517606 416820 517612 416832
rect 447928 416792 517612 416820
rect 447928 416780 447934 416792
rect 517606 416780 517612 416792
rect 517664 416780 517670 416832
rect 448974 415420 448980 415472
rect 449032 415460 449038 415472
rect 517514 415460 517520 415472
rect 449032 415432 517520 415460
rect 449032 415420 449038 415432
rect 517514 415420 517520 415432
rect 517572 415420 517578 415472
rect 449066 413992 449072 414044
rect 449124 414032 449130 414044
rect 517514 414032 517520 414044
rect 449124 414004 517520 414032
rect 449124 413992 449130 414004
rect 517514 413992 517520 414004
rect 517572 413992 517578 414044
rect 450354 412632 450360 412684
rect 450412 412672 450418 412684
rect 517514 412672 517520 412684
rect 450412 412644 517520 412672
rect 450412 412632 450418 412644
rect 517514 412632 517520 412644
rect 517572 412632 517578 412684
rect 450262 411272 450268 411324
rect 450320 411312 450326 411324
rect 517514 411312 517520 411324
rect 450320 411284 517520 411312
rect 450320 411272 450326 411284
rect 517514 411272 517520 411284
rect 517572 411272 517578 411324
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 43438 411244 43444 411256
rect 3384 411216 43444 411244
rect 3384 411204 3390 411216
rect 43438 411204 43444 411216
rect 43496 411204 43502 411256
rect 447686 409844 447692 409896
rect 447744 409884 447750 409896
rect 517514 409884 517520 409896
rect 447744 409856 517520 409884
rect 447744 409844 447750 409856
rect 517514 409844 517520 409856
rect 517572 409844 517578 409896
rect 450170 408484 450176 408536
rect 450228 408524 450234 408536
rect 517514 408524 517520 408536
rect 450228 408496 517520 408524
rect 450228 408484 450234 408496
rect 517514 408484 517520 408496
rect 517572 408484 517578 408536
rect 449986 407192 449992 407244
rect 450044 407232 450050 407244
rect 517514 407232 517520 407244
rect 450044 407204 517520 407232
rect 450044 407192 450050 407204
rect 517514 407192 517520 407204
rect 517572 407192 517578 407244
rect 450078 407124 450084 407176
rect 450136 407164 450142 407176
rect 517606 407164 517612 407176
rect 450136 407136 517612 407164
rect 450136 407124 450142 407136
rect 517606 407124 517612 407136
rect 517664 407124 517670 407176
rect 449894 405696 449900 405748
rect 449952 405736 449958 405748
rect 517514 405736 517520 405748
rect 449952 405708 517520 405736
rect 449952 405696 449958 405708
rect 517514 405696 517520 405708
rect 517572 405696 517578 405748
rect 562502 405628 562508 405680
rect 562560 405668 562566 405680
rect 580166 405668 580172 405680
rect 562560 405640 580172 405668
rect 562560 405628 562566 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 447778 404336 447784 404388
rect 447836 404376 447842 404388
rect 517514 404376 517520 404388
rect 447836 404348 517520 404376
rect 447836 404336 447842 404348
rect 517514 404336 517520 404348
rect 517572 404336 517578 404388
rect 449158 402976 449164 403028
rect 449216 403016 449222 403028
rect 517698 403016 517704 403028
rect 449216 402988 517704 403016
rect 449216 402976 449222 402988
rect 517698 402976 517704 402988
rect 517756 402976 517762 403028
rect 449342 401616 449348 401668
rect 449400 401656 449406 401668
rect 517698 401656 517704 401668
rect 449400 401628 517704 401656
rect 449400 401616 449406 401628
rect 517698 401616 517704 401628
rect 517756 401616 517762 401668
rect 449526 400256 449532 400308
rect 449584 400296 449590 400308
rect 517698 400296 517704 400308
rect 449584 400268 517704 400296
rect 449584 400256 449590 400268
rect 517698 400256 517704 400268
rect 517756 400256 517762 400308
rect 449250 400188 449256 400240
rect 449308 400228 449314 400240
rect 517790 400228 517796 400240
rect 449308 400200 517796 400228
rect 449308 400188 449314 400200
rect 517790 400188 517796 400200
rect 517848 400188 517854 400240
rect 449618 398828 449624 398880
rect 449676 398868 449682 398880
rect 517698 398868 517704 398880
rect 449676 398840 517704 398868
rect 449676 398828 449682 398840
rect 517698 398828 517704 398840
rect 517756 398828 517762 398880
rect 449434 397468 449440 397520
rect 449492 397508 449498 397520
rect 517698 397508 517704 397520
rect 449492 397480 517704 397508
rect 449492 397468 449498 397480
rect 517698 397468 517704 397480
rect 517756 397468 517762 397520
rect 449710 396040 449716 396092
rect 449768 396080 449774 396092
rect 517698 396080 517704 396092
rect 449768 396052 517704 396080
rect 449768 396040 449774 396052
rect 517698 396040 517704 396052
rect 517756 396040 517762 396092
rect 450814 394748 450820 394800
rect 450872 394788 450878 394800
rect 517698 394788 517704 394800
rect 450872 394760 517704 394788
rect 450872 394748 450878 394760
rect 517698 394748 517704 394760
rect 517756 394748 517762 394800
rect 449802 394680 449808 394732
rect 449860 394720 449866 394732
rect 517790 394720 517796 394732
rect 449860 394692 517796 394720
rect 449860 394680 449866 394692
rect 517790 394680 517796 394692
rect 517848 394680 517854 394732
rect 447042 393320 447048 393372
rect 447100 393360 447106 393372
rect 517698 393360 517704 393372
rect 447100 393332 517704 393360
rect 447100 393320 447106 393332
rect 517698 393320 517704 393332
rect 517756 393320 517762 393372
rect 448146 392096 448152 392148
rect 448204 392136 448210 392148
rect 517698 392136 517704 392148
rect 448204 392108 517704 392136
rect 448204 392096 448210 392108
rect 517698 392096 517704 392108
rect 517756 392096 517762 392148
rect 447962 392028 447968 392080
rect 448020 392068 448026 392080
rect 517882 392068 517888 392080
rect 448020 392040 517888 392068
rect 448020 392028 448026 392040
rect 517882 392028 517888 392040
rect 517940 392028 517946 392080
rect 446950 391960 446956 392012
rect 447008 392000 447014 392012
rect 517974 392000 517980 392012
rect 447008 391972 517980 392000
rect 447008 391960 447014 391972
rect 517974 391960 517980 391972
rect 518032 391960 518038 392012
rect 448054 390600 448060 390652
rect 448112 390640 448118 390652
rect 517698 390640 517704 390652
rect 448112 390612 517704 390640
rect 448112 390600 448118 390612
rect 517698 390600 517704 390612
rect 517756 390600 517762 390652
rect 446858 390532 446864 390584
rect 446916 390572 446922 390584
rect 517882 390572 517888 390584
rect 446916 390544 517888 390572
rect 446916 390532 446922 390544
rect 517882 390532 517888 390544
rect 517940 390532 517946 390584
rect 448238 389240 448244 389292
rect 448296 389280 448302 389292
rect 517698 389280 517704 389292
rect 448296 389252 517704 389280
rect 448296 389240 448302 389252
rect 517698 389240 517704 389252
rect 517756 389240 517762 389292
rect 446766 389172 446772 389224
rect 446824 389212 446830 389224
rect 517882 389212 517888 389224
rect 446824 389184 517888 389212
rect 446824 389172 446830 389184
rect 517882 389172 517888 389184
rect 517940 389172 517946 389224
rect 448330 387948 448336 388000
rect 448388 387988 448394 388000
rect 517882 387988 517888 388000
rect 448388 387960 517888 387988
rect 448388 387948 448394 387960
rect 517882 387948 517888 387960
rect 517940 387948 517946 388000
rect 446674 387880 446680 387932
rect 446732 387920 446738 387932
rect 517698 387920 517704 387932
rect 446732 387892 517704 387920
rect 446732 387880 446738 387892
rect 517698 387880 517704 387892
rect 517756 387880 517762 387932
rect 446582 387812 446588 387864
rect 446640 387852 446646 387864
rect 517974 387852 517980 387864
rect 446640 387824 517980 387852
rect 446640 387812 446646 387824
rect 517974 387812 517980 387824
rect 518032 387812 518038 387864
rect 448422 386452 448428 386504
rect 448480 386492 448486 386504
rect 517882 386492 517888 386504
rect 448480 386464 517888 386492
rect 448480 386452 448486 386464
rect 517882 386452 517888 386464
rect 517940 386452 517946 386504
rect 446490 386384 446496 386436
rect 446548 386424 446554 386436
rect 517698 386424 517704 386436
rect 446548 386396 517704 386424
rect 446548 386384 446554 386396
rect 517698 386384 517704 386396
rect 517756 386384 517762 386436
rect 517606 379856 517612 379908
rect 517664 379896 517670 379908
rect 550634 379896 550640 379908
rect 517664 379868 550640 379896
rect 517664 379856 517670 379868
rect 550634 379856 550640 379868
rect 550692 379856 550698 379908
rect 563882 379448 563888 379500
rect 563940 379488 563946 379500
rect 580166 379488 580172 379500
rect 563940 379460 580172 379488
rect 563940 379448 563946 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 519354 379108 519360 379160
rect 519412 379148 519418 379160
rect 549622 379148 549628 379160
rect 519412 379120 549628 379148
rect 519412 379108 519418 379120
rect 549622 379108 549628 379120
rect 549680 379108 549686 379160
rect 519078 379040 519084 379092
rect 519136 379080 519142 379092
rect 549714 379080 549720 379092
rect 519136 379052 549720 379080
rect 519136 379040 519142 379052
rect 549714 379040 549720 379052
rect 549772 379040 549778 379092
rect 518986 378972 518992 379024
rect 519044 379012 519050 379024
rect 549806 379012 549812 379024
rect 519044 378984 549812 379012
rect 519044 378972 519050 378984
rect 549806 378972 549812 378984
rect 549864 378972 549870 379024
rect 519446 378904 519452 378956
rect 519504 378944 519510 378956
rect 550726 378944 550732 378956
rect 519504 378916 550732 378944
rect 519504 378904 519510 378916
rect 550726 378904 550732 378916
rect 550784 378904 550790 378956
rect 519170 378836 519176 378888
rect 519228 378876 519234 378888
rect 550818 378876 550824 378888
rect 519228 378848 550824 378876
rect 519228 378836 519234 378848
rect 550818 378836 550824 378848
rect 550876 378836 550882 378888
rect 519262 378768 519268 378820
rect 519320 378808 519326 378820
rect 550910 378808 550916 378820
rect 519320 378780 550916 378808
rect 519320 378768 519326 378780
rect 550910 378768 550916 378780
rect 550968 378768 550974 378820
rect 521562 378020 521568 378072
rect 521620 378060 521626 378072
rect 523034 378060 523040 378072
rect 521620 378032 523040 378060
rect 521620 378020 521626 378032
rect 523034 378020 523040 378032
rect 523092 378020 523098 378072
rect 521286 377680 521292 377732
rect 521344 377720 521350 377732
rect 533338 377720 533344 377732
rect 521344 377692 533344 377720
rect 521344 377680 521350 377692
rect 533338 377680 533344 377692
rect 533396 377680 533402 377732
rect 524322 377612 524328 377664
rect 524380 377652 524386 377664
rect 549898 377652 549904 377664
rect 524380 377624 549904 377652
rect 524380 377612 524386 377624
rect 549898 377612 549904 377624
rect 549956 377612 549962 377664
rect 523402 377544 523408 377596
rect 523460 377584 523466 377596
rect 549990 377584 549996 377596
rect 523460 377556 549996 377584
rect 523460 377544 523466 377556
rect 549990 377544 549996 377556
rect 550048 377544 550054 377596
rect 524046 377476 524052 377528
rect 524104 377516 524110 377528
rect 551462 377516 551468 377528
rect 524104 377488 551468 377516
rect 524104 377476 524110 377488
rect 551462 377476 551468 377488
rect 551520 377476 551526 377528
rect 520366 377408 520372 377460
rect 520424 377448 520430 377460
rect 549254 377448 549260 377460
rect 520424 377420 549260 377448
rect 520424 377408 520430 377420
rect 549254 377408 549260 377420
rect 549312 377408 549318 377460
rect 524690 376116 524696 376168
rect 524748 376156 524754 376168
rect 550082 376156 550088 376168
rect 524748 376128 550088 376156
rect 524748 376116 524754 376128
rect 550082 376116 550088 376128
rect 550140 376116 550146 376168
rect 523126 376048 523132 376100
rect 523184 376088 523190 376100
rect 551278 376088 551284 376100
rect 523184 376060 551284 376088
rect 523184 376048 523190 376060
rect 551278 376048 551284 376060
rect 551336 376048 551342 376100
rect 523034 375980 523040 376032
rect 523092 376020 523098 376032
rect 552106 376020 552112 376032
rect 523092 375992 552112 376020
rect 523092 375980 523098 375992
rect 552106 375980 552112 375992
rect 552164 375980 552170 376032
rect 523770 374756 523776 374808
rect 523828 374796 523834 374808
rect 551370 374796 551376 374808
rect 523828 374768 551376 374796
rect 523828 374756 523834 374768
rect 551370 374756 551376 374768
rect 551428 374756 551434 374808
rect 520642 374688 520648 374740
rect 520700 374728 520706 374740
rect 551186 374728 551192 374740
rect 520700 374700 551192 374728
rect 520700 374688 520706 374700
rect 551186 374688 551192 374700
rect 551244 374688 551250 374740
rect 520090 374620 520096 374672
rect 520148 374660 520154 374672
rect 551094 374660 551100 374672
rect 520148 374632 551100 374660
rect 520148 374620 520154 374632
rect 551094 374620 551100 374632
rect 551152 374620 551158 374672
rect 533338 371900 533344 371952
rect 533396 371940 533402 371952
rect 552014 371940 552020 371952
rect 533396 371912 552020 371940
rect 533396 371900 533402 371912
rect 552014 371900 552020 371912
rect 552072 371900 552078 371952
rect 521010 371832 521016 371884
rect 521068 371872 521074 371884
rect 549346 371872 549352 371884
rect 521068 371844 549352 371872
rect 521068 371832 521074 371844
rect 549346 371832 549352 371844
rect 549404 371832 549410 371884
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 222194 371260 222200 371272
rect 3384 371232 222200 371260
rect 3384 371220 3390 371232
rect 222194 371220 222200 371232
rect 222252 371260 222258 371272
rect 223482 371260 223488 371272
rect 222252 371232 223488 371260
rect 222252 371220 222258 371232
rect 223482 371220 223488 371232
rect 223540 371220 223546 371272
rect 522850 371152 522856 371204
rect 522908 371192 522914 371204
rect 552474 371192 552480 371204
rect 522908 371164 552480 371192
rect 522908 371152 522914 371164
rect 552474 371152 552480 371164
rect 552532 371152 552538 371204
rect 522482 371084 522488 371136
rect 522540 371124 522546 371136
rect 552382 371124 552388 371136
rect 522540 371096 552388 371124
rect 522540 371084 522546 371096
rect 552382 371084 552388 371096
rect 552440 371084 552446 371136
rect 522206 371016 522212 371068
rect 522264 371056 522270 371068
rect 552290 371056 552296 371068
rect 522264 371028 552296 371056
rect 522264 371016 522270 371028
rect 552290 371016 552296 371028
rect 552348 371016 552354 371068
rect 521930 370948 521936 371000
rect 521988 370988 521994 371000
rect 552198 370988 552204 371000
rect 521988 370960 552204 370988
rect 521988 370948 521994 370960
rect 552198 370948 552204 370960
rect 552256 370948 552262 371000
rect 518894 370880 518900 370932
rect 518952 370920 518958 370932
rect 549530 370920 549536 370932
rect 518952 370892 549536 370920
rect 518952 370880 518958 370892
rect 549530 370880 549536 370892
rect 549588 370880 549594 370932
rect 517514 370812 517520 370864
rect 517572 370852 517578 370864
rect 549438 370852 549444 370864
rect 517572 370824 549444 370852
rect 517572 370812 517578 370824
rect 549438 370812 549444 370824
rect 549496 370812 549502 370864
rect 518250 370744 518256 370796
rect 518308 370784 518314 370796
rect 551002 370784 551008 370796
rect 518308 370756 551008 370784
rect 518308 370744 518314 370756
rect 551002 370744 551008 370756
rect 551060 370744 551066 370796
rect 518710 370676 518716 370728
rect 518768 370716 518774 370728
rect 553578 370716 553584 370728
rect 518768 370688 553584 370716
rect 518768 370676 518774 370688
rect 553578 370676 553584 370688
rect 553636 370676 553642 370728
rect 518802 370608 518808 370660
rect 518860 370648 518866 370660
rect 553670 370648 553676 370660
rect 518860 370620 553676 370648
rect 518860 370608 518866 370620
rect 553670 370608 553676 370620
rect 553728 370608 553734 370660
rect 514662 370540 514668 370592
rect 514720 370580 514726 370592
rect 553762 370580 553768 370592
rect 514720 370552 553768 370580
rect 514720 370540 514726 370552
rect 553762 370540 553768 370552
rect 553820 370540 553826 370592
rect 450722 370472 450728 370524
rect 450780 370512 450786 370524
rect 518158 370512 518164 370524
rect 450780 370484 518164 370512
rect 450780 370472 450786 370484
rect 518158 370472 518164 370484
rect 518216 370472 518222 370524
rect 518618 370472 518624 370524
rect 518676 370512 518682 370524
rect 553486 370512 553492 370524
rect 518676 370484 553492 370512
rect 518676 370472 518682 370484
rect 553486 370472 553492 370484
rect 553544 370472 553550 370524
rect 3050 358708 3056 358760
rect 3108 358748 3114 358760
rect 87598 358748 87604 358760
rect 3108 358720 87604 358748
rect 3108 358708 3114 358720
rect 87598 358708 87604 358720
rect 87656 358708 87662 358760
rect 560754 353200 560760 353252
rect 560812 353240 560818 353252
rect 579614 353240 579620 353252
rect 560812 353212 579620 353240
rect 560812 353200 560818 353212
rect 579614 353200 579620 353212
rect 579672 353200 579678 353252
rect 549898 352520 549904 352572
rect 549956 352560 549962 352572
rect 560754 352560 560760 352572
rect 549956 352532 560760 352560
rect 549956 352520 549962 352532
rect 560754 352520 560760 352532
rect 560812 352520 560818 352572
rect 2958 346332 2964 346384
rect 3016 346372 3022 346384
rect 444742 346372 444748 346384
rect 3016 346344 444748 346372
rect 3016 346332 3022 346344
rect 444742 346332 444748 346344
rect 444800 346332 444806 346384
rect 563790 325592 563796 325644
rect 563848 325632 563854 325644
rect 580166 325632 580172 325644
rect 563848 325604 580172 325632
rect 563848 325592 563854 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 226334 320084 226340 320136
rect 226392 320124 226398 320136
rect 226978 320124 226984 320136
rect 226392 320096 226984 320124
rect 226392 320084 226398 320096
rect 226978 320084 226984 320096
rect 227036 320084 227042 320136
rect 3326 319404 3332 319456
rect 3384 319444 3390 319456
rect 226334 319444 226340 319456
rect 3384 319416 226340 319444
rect 3384 319404 3390 319416
rect 226334 319404 226340 319416
rect 226392 319404 226398 319456
rect 566458 313216 566464 313268
rect 566516 313256 566522 313268
rect 580166 313256 580172 313268
rect 566516 313228 580172 313256
rect 566516 313216 566522 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 175918 306320 175924 306332
rect 3384 306292 175924 306320
rect 3384 306280 3390 306292
rect 175918 306280 175924 306292
rect 175976 306280 175982 306332
rect 561582 299412 561588 299464
rect 561640 299452 561646 299464
rect 580166 299452 580172 299464
rect 561640 299424 580172 299452
rect 561640 299412 561646 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 113174 298732 113180 298784
rect 113232 298772 113238 298784
rect 560662 298772 560668 298784
rect 113232 298744 560668 298772
rect 113232 298732 113238 298744
rect 560662 298732 560668 298744
rect 560720 298772 560726 298784
rect 561582 298772 561588 298784
rect 560720 298744 561588 298772
rect 560720 298732 560726 298744
rect 561582 298732 561588 298744
rect 561640 298732 561646 298784
rect 446490 298052 446496 298104
rect 446548 298092 446554 298104
rect 460750 298092 460756 298104
rect 446548 298064 460756 298092
rect 446548 298052 446554 298064
rect 460750 298052 460756 298064
rect 460808 298052 460814 298104
rect 545206 298052 545212 298104
rect 545264 298092 545270 298104
rect 553394 298092 553400 298104
rect 545264 298064 553400 298092
rect 545264 298052 545270 298064
rect 553394 298052 553400 298064
rect 553452 298052 553458 298104
rect 450814 297984 450820 298036
rect 450872 298024 450878 298036
rect 482646 298024 482652 298036
rect 450872 297996 482652 298024
rect 450872 297984 450878 297996
rect 482646 297984 482652 297996
rect 482704 297984 482710 298036
rect 535822 297984 535828 298036
rect 535880 298024 535886 298036
rect 553486 298024 553492 298036
rect 535880 297996 553492 298024
rect 535880 297984 535886 297996
rect 553486 297984 553492 297996
rect 553544 297984 553550 298036
rect 446950 297916 446956 297968
rect 447008 297956 447014 297968
rect 476390 297956 476396 297968
rect 447008 297928 476396 297956
rect 447008 297916 447014 297928
rect 476390 297916 476396 297928
rect 476448 297916 476454 297968
rect 538950 297916 538956 297968
rect 539008 297956 539014 297968
rect 553578 297956 553584 297968
rect 539008 297928 553584 297956
rect 539008 297916 539014 297928
rect 553578 297916 553584 297928
rect 553636 297916 553642 297968
rect 446858 297848 446864 297900
rect 446916 297888 446922 297900
rect 473262 297888 473268 297900
rect 446916 297860 473268 297888
rect 446916 297848 446922 297860
rect 473262 297848 473268 297860
rect 473320 297848 473326 297900
rect 542078 297848 542084 297900
rect 542136 297888 542142 297900
rect 553670 297888 553676 297900
rect 542136 297860 553676 297888
rect 542136 297848 542142 297860
rect 553670 297848 553676 297860
rect 553728 297848 553734 297900
rect 446766 297780 446772 297832
rect 446824 297820 446830 297832
rect 470134 297820 470140 297832
rect 446824 297792 470140 297820
rect 446824 297780 446830 297792
rect 470134 297780 470140 297792
rect 470192 297780 470198 297832
rect 510798 297780 510804 297832
rect 510856 297820 510862 297832
rect 550910 297820 550916 297832
rect 510856 297792 550916 297820
rect 510856 297780 510862 297792
rect 550910 297780 550916 297792
rect 550968 297780 550974 297832
rect 446582 297712 446588 297764
rect 446640 297752 446646 297764
rect 467006 297752 467012 297764
rect 446640 297724 467012 297752
rect 446640 297712 446646 297724
rect 467006 297712 467012 297724
rect 467064 297712 467070 297764
rect 513926 297712 513932 297764
rect 513984 297752 513990 297764
rect 549806 297752 549812 297764
rect 513984 297724 549812 297752
rect 513984 297712 513990 297724
rect 549806 297712 549812 297724
rect 549864 297712 549870 297764
rect 446674 297644 446680 297696
rect 446732 297684 446738 297696
rect 463878 297684 463884 297696
rect 446732 297656 463884 297684
rect 446732 297644 446738 297656
rect 463878 297644 463884 297656
rect 463936 297644 463942 297696
rect 517054 297644 517060 297696
rect 517112 297684 517118 297696
rect 550634 297684 550640 297696
rect 517112 297656 550640 297684
rect 517112 297644 517118 297656
rect 550634 297644 550640 297656
rect 550692 297644 550698 297696
rect 447042 297576 447048 297628
rect 447100 297616 447106 297628
rect 479518 297616 479524 297628
rect 447100 297588 479524 297616
rect 447100 297576 447106 297588
rect 479518 297576 479524 297588
rect 479576 297576 479582 297628
rect 520182 297576 520188 297628
rect 520240 297616 520246 297628
rect 549530 297616 549536 297628
rect 520240 297588 549536 297616
rect 520240 297576 520246 297588
rect 549530 297576 549536 297588
rect 549588 297576 549594 297628
rect 523310 297508 523316 297560
rect 523368 297548 523374 297560
rect 551002 297548 551008 297560
rect 523368 297520 551008 297548
rect 523368 297508 523374 297520
rect 551002 297508 551008 297520
rect 551060 297508 551066 297560
rect 498286 297440 498292 297492
rect 498344 297480 498350 297492
rect 550726 297480 550732 297492
rect 498344 297452 550732 297480
rect 498344 297440 498350 297452
rect 550726 297440 550732 297452
rect 550784 297440 550790 297492
rect 501414 297372 501420 297424
rect 501472 297412 501478 297424
rect 549622 297412 549628 297424
rect 501472 297384 549628 297412
rect 501472 297372 501478 297384
rect 549622 297372 549628 297384
rect 549680 297372 549686 297424
rect 504542 297304 504548 297356
rect 504600 297344 504606 297356
rect 550818 297344 550824 297356
rect 504600 297316 550824 297344
rect 504600 297304 504606 297316
rect 550818 297304 550824 297316
rect 550876 297304 550882 297356
rect 507670 297236 507676 297288
rect 507728 297276 507734 297288
rect 549714 297276 549720 297288
rect 507728 297248 549720 297276
rect 507728 297236 507734 297248
rect 549714 297236 549720 297248
rect 549772 297236 549778 297288
rect 526438 297168 526444 297220
rect 526496 297208 526502 297220
rect 549438 297208 549444 297220
rect 526496 297180 549444 297208
rect 526496 297168 526502 297180
rect 549438 297168 549444 297180
rect 549496 297168 549502 297220
rect 3234 293904 3240 293956
rect 3292 293944 3298 293956
rect 444926 293944 444932 293956
rect 3292 293916 444932 293944
rect 3292 293904 3298 293916
rect 444926 293904 444932 293916
rect 444984 293904 444990 293956
rect 562410 273164 562416 273216
rect 562468 273204 562474 273216
rect 580166 273204 580172 273216
rect 562468 273176 580172 273204
rect 562468 273164 562474 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 231854 267180 231860 267232
rect 231912 267220 231918 267232
rect 232498 267220 232504 267232
rect 231912 267192 232504 267220
rect 231912 267180 231918 267192
rect 232498 267180 232504 267192
rect 232556 267180 232562 267232
rect 3326 266976 3332 267028
rect 3384 267016 3390 267028
rect 231854 267016 231860 267028
rect 3384 266988 231860 267016
rect 3384 266976 3390 266988
rect 231854 266976 231860 266988
rect 231912 266976 231918 267028
rect 563698 259360 563704 259412
rect 563756 259400 563762 259412
rect 579798 259400 579804 259412
rect 563756 259372 579804 259400
rect 563756 259360 563762 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 2958 255212 2964 255264
rect 3016 255252 3022 255264
rect 352558 255252 352564 255264
rect 3016 255224 352564 255252
rect 3016 255212 3022 255224
rect 352558 255212 352564 255224
rect 352616 255212 352622 255264
rect 560570 245556 560576 245608
rect 560628 245596 560634 245608
rect 580166 245596 580172 245608
rect 560628 245568 580172 245596
rect 560628 245556 560634 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 440878 244876 440884 244928
rect 440936 244916 440942 244928
rect 560570 244916 560576 244928
rect 440936 244888 560576 244916
rect 440936 244876 440942 244888
rect 560570 244876 560576 244888
rect 560628 244876 560634 244928
rect 109034 224204 109040 224256
rect 109092 224244 109098 224256
rect 440878 224244 440884 224256
rect 109092 224216 440884 224244
rect 109092 224204 109098 224216
rect 440878 224204 440884 224216
rect 440936 224204 440942 224256
rect 3326 214548 3332 214600
rect 3384 214588 3390 214600
rect 235994 214588 236000 214600
rect 3384 214560 236000 214588
rect 3384 214548 3390 214560
rect 235994 214548 236000 214560
rect 236052 214588 236058 214600
rect 236638 214588 236644 214600
rect 236052 214560 236644 214588
rect 236052 214548 236058 214560
rect 236638 214548 236644 214560
rect 236696 214548 236702 214600
rect 560478 206932 560484 206984
rect 560536 206972 560542 206984
rect 579798 206972 579804 206984
rect 560536 206944 579804 206972
rect 560536 206932 560542 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 103974 206252 103980 206304
rect 104032 206292 104038 206304
rect 560478 206292 560484 206304
rect 104032 206264 560484 206292
rect 104032 206252 104038 206264
rect 560478 206252 560484 206264
rect 560536 206252 560542 206304
rect 170306 203736 170312 203788
rect 170364 203776 170370 203788
rect 300118 203776 300124 203788
rect 170364 203748 300124 203776
rect 170364 203736 170370 203748
rect 300118 203736 300124 203748
rect 300176 203736 300182 203788
rect 40034 203668 40040 203720
rect 40092 203708 40098 203720
rect 189074 203708 189080 203720
rect 40092 203680 189080 203708
rect 40092 203668 40098 203680
rect 189074 203668 189080 203680
rect 189132 203668 189138 203720
rect 165614 203600 165620 203652
rect 165672 203640 165678 203652
rect 364978 203640 364984 203652
rect 165672 203612 364984 203640
rect 165672 203600 165678 203612
rect 364978 203600 364984 203612
rect 365036 203600 365042 203652
rect 4890 203532 4896 203584
rect 4948 203572 4954 203584
rect 218146 203572 218152 203584
rect 4948 203544 218152 203572
rect 4948 203532 4954 203544
rect 218146 203532 218152 203544
rect 218204 203532 218210 203584
rect 189074 202784 189080 202836
rect 189132 202824 189138 202836
rect 189718 202824 189724 202836
rect 189132 202796 189724 202824
rect 189132 202784 189138 202796
rect 189718 202784 189724 202796
rect 189776 202824 189782 202836
rect 445386 202824 445392 202836
rect 189776 202796 445392 202824
rect 189776 202784 189782 202796
rect 445386 202784 445392 202796
rect 445444 202784 445450 202836
rect 123662 202512 123668 202564
rect 123720 202552 123726 202564
rect 284938 202552 284944 202564
rect 123720 202524 284944 202552
rect 123720 202512 123726 202524
rect 284938 202512 284944 202524
rect 284996 202512 285002 202564
rect 156874 202444 156880 202496
rect 156932 202484 156938 202496
rect 445018 202484 445024 202496
rect 156932 202456 445024 202484
rect 156932 202444 156938 202456
rect 445018 202444 445024 202456
rect 445076 202444 445082 202496
rect 152090 202376 152096 202428
rect 152148 202416 152154 202428
rect 445110 202416 445116 202428
rect 152148 202388 445116 202416
rect 152148 202376 152154 202388
rect 445110 202376 445116 202388
rect 445168 202376 445174 202428
rect 147398 202308 147404 202360
rect 147456 202348 147462 202360
rect 445202 202348 445208 202360
rect 147456 202320 445208 202348
rect 147456 202308 147462 202320
rect 445202 202308 445208 202320
rect 445260 202308 445266 202360
rect 142614 202240 142620 202292
rect 142672 202280 142678 202292
rect 445294 202280 445300 202292
rect 142672 202252 445300 202280
rect 142672 202240 142678 202252
rect 445294 202240 445300 202252
rect 445352 202240 445358 202292
rect 175826 202172 175832 202224
rect 175884 202212 175890 202224
rect 235258 202212 235264 202224
rect 175884 202184 235264 202212
rect 175884 202172 175890 202184
rect 235258 202172 235264 202184
rect 235316 202172 235322 202224
rect 256050 202172 256056 202224
rect 256108 202212 256114 202224
rect 559926 202212 559932 202224
rect 256108 202184 559932 202212
rect 256108 202172 256114 202184
rect 559926 202172 559932 202184
rect 559984 202172 559990 202224
rect 118970 202104 118976 202156
rect 119028 202144 119034 202156
rect 549898 202144 549904 202156
rect 119028 202116 549904 202144
rect 119028 202104 119034 202116
rect 549898 202104 549904 202116
rect 549956 202104 549962 202156
rect 100018 201628 100024 201680
rect 100076 201668 100082 201680
rect 261570 201668 261576 201680
rect 100076 201640 261576 201668
rect 100076 201628 100082 201640
rect 261570 201628 261576 201640
rect 261628 201628 261634 201680
rect 95142 201560 95148 201612
rect 95200 201600 95206 201612
rect 260098 201600 260104 201612
rect 95200 201572 260104 201600
rect 95200 201560 95206 201572
rect 260098 201560 260104 201572
rect 260156 201560 260162 201612
rect 3786 201492 3792 201544
rect 3844 201532 3850 201544
rect 256050 201532 256056 201544
rect 3844 201504 256056 201532
rect 3844 201492 3850 201504
rect 256050 201492 256056 201504
rect 256108 201492 256114 201544
rect 561306 201424 561312 201476
rect 561364 201464 561370 201476
rect 564434 201464 564440 201476
rect 561364 201436 564440 201464
rect 561364 201424 561370 201436
rect 564434 201424 564440 201436
rect 564492 201424 564498 201476
rect 251358 200880 251364 200932
rect 251416 200920 251422 200932
rect 445570 200920 445576 200932
rect 251416 200892 445576 200920
rect 251416 200880 251422 200892
rect 445570 200880 445576 200892
rect 445628 200880 445634 200932
rect 246574 200812 246580 200864
rect 246632 200852 246638 200864
rect 445662 200852 445668 200864
rect 246632 200824 445668 200852
rect 246632 200812 246638 200824
rect 445662 200812 445668 200824
rect 445720 200812 445726 200864
rect 241882 200744 241888 200796
rect 241940 200784 241946 200796
rect 445478 200784 445484 200796
rect 241940 200756 445484 200784
rect 241940 200744 241946 200756
rect 445478 200744 445484 200756
rect 445536 200744 445542 200796
rect 85482 200472 85488 200524
rect 85540 200512 85546 200524
rect 261478 200512 261484 200524
rect 85540 200484 261484 200512
rect 85540 200472 85546 200484
rect 261478 200472 261484 200484
rect 261536 200472 261542 200524
rect 4890 200404 4896 200456
rect 4948 200444 4954 200456
rect 241882 200444 241888 200456
rect 4948 200416 241888 200444
rect 4948 200404 4954 200416
rect 241882 200404 241888 200416
rect 241940 200404 241946 200456
rect 3878 200336 3884 200388
rect 3936 200376 3942 200388
rect 246574 200376 246580 200388
rect 3936 200348 246580 200376
rect 3936 200336 3942 200348
rect 246574 200336 246580 200348
rect 246632 200336 246638 200388
rect 3694 200268 3700 200320
rect 3752 200308 3758 200320
rect 251358 200308 251364 200320
rect 3752 200280 251364 200308
rect 3752 200268 3758 200280
rect 251358 200268 251364 200280
rect 251416 200268 251422 200320
rect 90542 200200 90548 200252
rect 90600 200240 90606 200252
rect 438118 200240 438124 200252
rect 90600 200212 438124 200240
rect 90600 200200 90606 200212
rect 438118 200200 438124 200212
rect 438176 200200 438182 200252
rect 81066 200132 81072 200184
rect 81124 200172 81130 200184
rect 561306 200172 561312 200184
rect 81124 200144 561312 200172
rect 81124 200132 81130 200144
rect 561306 200132 561312 200144
rect 561364 200132 561370 200184
rect 562318 193128 562324 193180
rect 562376 193168 562382 193180
rect 579614 193168 579620 193180
rect 562376 193140 579620 193168
rect 562376 193128 562382 193140
rect 579614 193128 579620 193140
rect 579672 193128 579678 193180
rect 569218 179324 569224 179376
rect 569276 179364 569282 179376
rect 579614 179364 579620 179376
rect 569276 179336 579620 179364
rect 569276 179324 569282 179336
rect 579614 179324 579620 179336
rect 579672 179324 579678 179376
rect 261570 166948 261576 167000
rect 261628 166988 261634 167000
rect 560386 166988 560392 167000
rect 261628 166960 560392 166988
rect 261628 166948 261634 166960
rect 560386 166948 560392 166960
rect 560444 166988 560450 167000
rect 580166 166988 580172 167000
rect 560444 166960 580172 166988
rect 560444 166948 560450 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 2774 162936 2780 162988
rect 2832 162976 2838 162988
rect 4890 162976 4896 162988
rect 2832 162948 4896 162976
rect 2832 162936 2838 162948
rect 4890 162936 4896 162948
rect 4948 162936 4954 162988
rect 2774 150152 2780 150204
rect 2832 150192 2838 150204
rect 4982 150192 4988 150204
rect 2832 150164 4988 150192
rect 2832 150152 2838 150164
rect 4982 150152 4988 150164
rect 5040 150152 5046 150204
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 79318 137952 79324 137964
rect 3568 137924 79324 137952
rect 3568 137912 3574 137924
rect 79318 137912 79324 137924
rect 79376 137912 79382 137964
rect 260098 126896 260104 126948
rect 260156 126936 260162 126948
rect 560018 126936 560024 126948
rect 260156 126908 560024 126936
rect 260156 126896 260162 126908
rect 560018 126896 560024 126908
rect 560076 126936 560082 126948
rect 580166 126936 580172 126948
rect 560076 126908 580172 126936
rect 560076 126896 560082 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 561214 113092 561220 113144
rect 561272 113132 561278 113144
rect 579614 113132 579620 113144
rect 561272 113104 579620 113132
rect 561272 113092 561278 113104
rect 579614 113092 579620 113104
rect 579672 113092 579678 113144
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 438118 86912 438124 86964
rect 438176 86952 438182 86964
rect 580166 86952 580172 86964
rect 438176 86924 547874 86952
rect 438176 86912 438182 86924
rect 547846 86884 547874 86924
rect 567166 86924 580172 86952
rect 560294 86884 560300 86896
rect 547846 86856 560300 86884
rect 560294 86844 560300 86856
rect 560352 86884 560358 86896
rect 567166 86884 567194 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 560352 86856 567194 86884
rect 560352 86844 560358 86856
rect 2958 85484 2964 85536
rect 3016 85524 3022 85536
rect 77938 85524 77944 85536
rect 3016 85496 77944 85524
rect 3016 85484 3022 85496
rect 77938 85484 77944 85496
rect 77996 85484 78002 85536
rect 80744 79880 80750 79892
rect 80072 79852 80750 79880
rect 80072 79824 80100 79852
rect 80744 79840 80750 79852
rect 80802 79840 80808 79892
rect 89806 79840 89812 79892
rect 89864 79880 89870 79892
rect 90680 79880 90686 79892
rect 89864 79852 90686 79880
rect 89864 79840 89870 79852
rect 90680 79840 90686 79852
rect 90738 79840 90744 79892
rect 96706 79840 96712 79892
rect 96764 79880 96770 79892
rect 97580 79880 97586 79892
rect 96764 79852 97586 79880
rect 96764 79840 96770 79852
rect 97580 79840 97586 79852
rect 97638 79840 97644 79892
rect 98086 79840 98092 79892
rect 98144 79880 98150 79892
rect 99052 79880 99058 79892
rect 98144 79852 99058 79880
rect 98144 79840 98150 79852
rect 99052 79840 99058 79852
rect 99110 79840 99116 79892
rect 121546 79840 121552 79892
rect 121604 79880 121610 79892
rect 122420 79880 122426 79892
rect 121604 79852 122426 79880
rect 121604 79840 121610 79852
rect 122420 79840 122426 79852
rect 122478 79840 122484 79892
rect 123524 79840 123530 79892
rect 123582 79840 123588 79892
rect 139992 79880 139998 79892
rect 139596 79852 139998 79880
rect 80054 79772 80060 79824
rect 80112 79772 80118 79824
rect 80146 79772 80152 79824
rect 80204 79812 80210 79824
rect 81112 79812 81118 79824
rect 80204 79784 81118 79812
rect 80204 79772 80210 79784
rect 81112 79772 81118 79784
rect 81170 79772 81176 79824
rect 81618 79772 81624 79824
rect 81676 79812 81682 79824
rect 82216 79812 82222 79824
rect 81676 79784 82222 79812
rect 81676 79772 81682 79784
rect 82216 79772 82222 79784
rect 82274 79772 82280 79824
rect 89714 79772 89720 79824
rect 89772 79812 89778 79824
rect 90312 79812 90318 79824
rect 89772 79784 90318 79812
rect 89772 79772 89778 79784
rect 90312 79772 90318 79784
rect 90370 79772 90376 79824
rect 96614 79772 96620 79824
rect 96672 79812 96678 79824
rect 97212 79812 97218 79824
rect 96672 79784 97218 79812
rect 96672 79772 96678 79784
rect 97212 79772 97218 79784
rect 97270 79772 97276 79824
rect 98178 79772 98184 79824
rect 98236 79812 98242 79824
rect 98684 79812 98690 79824
rect 98236 79784 98690 79812
rect 98236 79772 98242 79784
rect 98684 79772 98690 79784
rect 98742 79772 98748 79824
rect 99558 79772 99564 79824
rect 99616 79812 99622 79824
rect 100524 79812 100530 79824
rect 99616 79784 100530 79812
rect 99616 79772 99622 79784
rect 100524 79772 100530 79784
rect 100582 79772 100588 79824
rect 103606 79772 103612 79824
rect 103664 79812 103670 79824
rect 104480 79812 104486 79824
rect 103664 79784 104486 79812
rect 103664 79772 103670 79784
rect 104480 79772 104486 79784
rect 104538 79772 104544 79824
rect 106366 79772 106372 79824
rect 106424 79812 106430 79824
rect 107056 79812 107062 79824
rect 106424 79784 107062 79812
rect 106424 79772 106430 79784
rect 107056 79772 107062 79784
rect 107114 79772 107120 79824
rect 111978 79772 111984 79824
rect 112036 79812 112042 79824
rect 112576 79812 112582 79824
rect 112036 79784 112582 79812
rect 112036 79772 112042 79784
rect 112576 79772 112582 79784
rect 112634 79772 112640 79824
rect 116026 79772 116032 79824
rect 116084 79812 116090 79824
rect 116900 79812 116906 79824
rect 116084 79784 116906 79812
rect 116084 79772 116090 79784
rect 116900 79772 116906 79784
rect 116958 79772 116964 79824
rect 121454 79772 121460 79824
rect 121512 79812 121518 79824
rect 122052 79812 122058 79824
rect 121512 79784 122058 79812
rect 121512 79772 121518 79784
rect 122052 79772 122058 79784
rect 122110 79772 122116 79824
rect 79962 79636 79968 79688
rect 80020 79676 80026 79688
rect 80238 79676 80244 79688
rect 80020 79648 80244 79676
rect 80020 79636 80026 79648
rect 80238 79636 80244 79648
rect 80296 79636 80302 79688
rect 122834 79636 122840 79688
rect 122892 79676 122898 79688
rect 123542 79676 123570 79840
rect 139596 79824 139624 79852
rect 139992 79840 139998 79852
rect 140050 79840 140056 79892
rect 146294 79840 146300 79892
rect 146352 79880 146358 79892
rect 147260 79880 147266 79892
rect 146352 79852 147266 79880
rect 146352 79840 146358 79852
rect 147260 79840 147266 79852
rect 147318 79840 147324 79892
rect 151814 79840 151820 79892
rect 151872 79880 151878 79892
rect 152688 79880 152694 79892
rect 151872 79852 152694 79880
rect 151872 79840 151878 79852
rect 152688 79840 152694 79852
rect 152746 79840 152752 79892
rect 157334 79840 157340 79892
rect 157392 79880 157398 79892
rect 157840 79880 157846 79892
rect 157392 79852 157846 79880
rect 157392 79840 157398 79852
rect 157840 79840 157846 79852
rect 157898 79840 157904 79892
rect 158208 79840 158214 79892
rect 158266 79840 158272 79892
rect 170628 79880 170634 79892
rect 169864 79852 170634 79880
rect 124306 79772 124312 79824
rect 124364 79812 124370 79824
rect 125364 79812 125370 79824
rect 124364 79784 125370 79812
rect 124364 79772 124370 79784
rect 125364 79772 125370 79784
rect 125422 79772 125428 79824
rect 126974 79772 126980 79824
rect 127032 79812 127038 79824
rect 128216 79812 128222 79824
rect 127032 79784 128222 79812
rect 127032 79772 127038 79784
rect 128216 79772 128222 79784
rect 128274 79772 128280 79824
rect 129918 79772 129924 79824
rect 129976 79812 129982 79824
rect 130792 79812 130798 79824
rect 129976 79784 130798 79812
rect 129976 79772 129982 79784
rect 130792 79772 130798 79784
rect 130850 79772 130856 79824
rect 132494 79772 132500 79824
rect 132552 79812 132558 79824
rect 133000 79812 133006 79824
rect 132552 79784 133006 79812
rect 132552 79772 132558 79784
rect 133000 79772 133006 79784
rect 133058 79772 133064 79824
rect 133966 79772 133972 79824
rect 134024 79812 134030 79824
rect 134840 79812 134846 79824
rect 134024 79784 134846 79812
rect 134024 79772 134030 79784
rect 134840 79772 134846 79784
rect 134898 79772 134904 79824
rect 139578 79772 139584 79824
rect 139636 79772 139642 79824
rect 140774 79772 140780 79824
rect 140832 79812 140838 79824
rect 141740 79812 141746 79824
rect 140832 79784 141746 79812
rect 140832 79772 140838 79784
rect 141740 79772 141746 79784
rect 141798 79772 141804 79824
rect 144914 79772 144920 79824
rect 144972 79812 144978 79824
rect 146156 79812 146162 79824
rect 144972 79784 146162 79812
rect 144972 79772 144978 79784
rect 146156 79772 146162 79784
rect 146214 79772 146220 79824
rect 146386 79772 146392 79824
rect 146444 79812 146450 79824
rect 146892 79812 146898 79824
rect 146444 79784 146898 79812
rect 146444 79772 146450 79784
rect 146892 79772 146898 79784
rect 146950 79772 146956 79824
rect 147858 79772 147864 79824
rect 147916 79812 147922 79824
rect 148732 79812 148738 79824
rect 147916 79784 148738 79812
rect 147916 79772 147922 79784
rect 148732 79772 148738 79784
rect 148790 79772 148796 79824
rect 151998 79772 152004 79824
rect 152056 79812 152062 79824
rect 153056 79812 153062 79824
rect 152056 79784 153062 79812
rect 152056 79772 152062 79784
rect 153056 79772 153062 79784
rect 153114 79772 153120 79824
rect 153194 79772 153200 79824
rect 153252 79812 153258 79824
rect 154160 79812 154166 79824
rect 153252 79784 154166 79812
rect 153252 79772 153258 79784
rect 154160 79772 154166 79784
rect 154218 79772 154224 79824
rect 156138 79772 156144 79824
rect 156196 79812 156202 79824
rect 157104 79812 157110 79824
rect 156196 79784 157110 79812
rect 156196 79772 156202 79784
rect 157104 79772 157110 79784
rect 157162 79772 157168 79824
rect 122892 79648 123570 79676
rect 122892 79636 122898 79648
rect 157426 79636 157432 79688
rect 157484 79676 157490 79688
rect 158226 79676 158254 79840
rect 169864 79824 169892 79852
rect 170628 79840 170634 79852
rect 170686 79840 170692 79892
rect 174308 79880 174314 79892
rect 173912 79852 174314 79880
rect 162854 79772 162860 79824
rect 162912 79812 162918 79824
rect 163728 79812 163734 79824
rect 162912 79784 163734 79812
rect 162912 79772 162918 79784
rect 163728 79772 163734 79784
rect 163786 79772 163792 79824
rect 164234 79772 164240 79824
rect 164292 79812 164298 79824
rect 164740 79812 164746 79824
rect 164292 79784 164746 79812
rect 164292 79772 164298 79784
rect 164740 79772 164746 79784
rect 164798 79772 164804 79824
rect 166994 79772 167000 79824
rect 167052 79812 167058 79824
rect 168052 79812 168058 79824
rect 167052 79784 168058 79812
rect 167052 79772 167058 79784
rect 168052 79772 168058 79784
rect 168110 79772 168116 79824
rect 169846 79772 169852 79824
rect 169904 79772 169910 79824
rect 171226 79772 171232 79824
rect 171284 79812 171290 79824
rect 172100 79812 172106 79824
rect 171284 79784 172106 79812
rect 171284 79772 171290 79784
rect 172100 79772 172106 79784
rect 172158 79772 172164 79824
rect 173912 79688 173940 79852
rect 174308 79840 174314 79852
rect 174366 79840 174372 79892
rect 174676 79840 174682 79892
rect 174734 79840 174740 79892
rect 183646 79840 183652 79892
rect 183704 79880 183710 79892
rect 184520 79880 184526 79892
rect 183704 79852 184526 79880
rect 183704 79840 183710 79852
rect 184520 79840 184526 79852
rect 184578 79840 184584 79892
rect 189074 79840 189080 79892
rect 189132 79880 189138 79892
rect 189948 79880 189954 79892
rect 189132 79852 189954 79880
rect 189132 79840 189138 79852
rect 189948 79840 189954 79852
rect 190006 79840 190012 79892
rect 200528 79840 200534 79892
rect 200586 79840 200592 79892
rect 200896 79840 200902 79892
rect 200954 79840 200960 79892
rect 206416 79840 206422 79892
rect 206474 79840 206480 79892
rect 225368 79880 225374 79892
rect 224972 79852 225374 79880
rect 157484 79648 158254 79676
rect 157484 79636 157490 79648
rect 173894 79636 173900 79688
rect 173952 79636 173958 79688
rect 173986 79636 173992 79688
rect 174044 79676 174050 79688
rect 174694 79676 174722 79840
rect 176654 79772 176660 79824
rect 176712 79812 176718 79824
rect 177528 79812 177534 79824
rect 176712 79784 177534 79812
rect 176712 79772 176718 79784
rect 177528 79772 177534 79784
rect 177586 79772 177592 79824
rect 178034 79772 178040 79824
rect 178092 79812 178098 79824
rect 178632 79812 178638 79824
rect 178092 79784 178638 79812
rect 178092 79772 178098 79784
rect 178632 79772 178638 79784
rect 178690 79772 178696 79824
rect 182174 79772 182180 79824
rect 182232 79812 182238 79824
rect 183048 79812 183054 79824
rect 182232 79784 183054 79812
rect 182232 79772 182238 79784
rect 183048 79772 183054 79784
rect 183106 79772 183112 79824
rect 183554 79772 183560 79824
rect 183612 79812 183618 79824
rect 184152 79812 184158 79824
rect 183612 79784 184158 79812
rect 183612 79772 183618 79784
rect 184152 79772 184158 79784
rect 184210 79772 184216 79824
rect 187786 79772 187792 79824
rect 187844 79812 187850 79824
rect 188844 79812 188850 79824
rect 187844 79784 188850 79812
rect 187844 79772 187850 79784
rect 188844 79772 188850 79784
rect 188902 79772 188908 79824
rect 190454 79772 190460 79824
rect 190512 79812 190518 79824
rect 191052 79812 191058 79824
rect 190512 79784 191058 79812
rect 190512 79772 190518 79784
rect 191052 79772 191058 79784
rect 191110 79772 191116 79824
rect 193398 79772 193404 79824
rect 193456 79812 193462 79824
rect 194364 79812 194370 79824
rect 193456 79784 194370 79812
rect 193456 79772 193462 79784
rect 194364 79772 194370 79784
rect 194422 79772 194428 79824
rect 194594 79772 194600 79824
rect 194652 79812 194658 79824
rect 195468 79812 195474 79824
rect 194652 79784 195474 79812
rect 194652 79772 194658 79784
rect 195468 79772 195474 79784
rect 195526 79772 195532 79824
rect 198918 79772 198924 79824
rect 198976 79812 198982 79824
rect 199884 79812 199890 79824
rect 198976 79784 199890 79812
rect 198976 79772 198982 79784
rect 199884 79772 199890 79784
rect 199942 79772 199948 79824
rect 200546 79744 200574 79840
rect 200132 79716 200574 79744
rect 200132 79688 200160 79716
rect 174044 79648 174722 79676
rect 174044 79636 174050 79648
rect 200114 79636 200120 79688
rect 200172 79636 200178 79688
rect 200206 79636 200212 79688
rect 200264 79676 200270 79688
rect 200914 79676 200942 79840
rect 204346 79772 204352 79824
rect 204404 79812 204410 79824
rect 205312 79812 205318 79824
rect 204404 79784 205318 79812
rect 204404 79772 204410 79784
rect 205312 79772 205318 79784
rect 205370 79772 205376 79824
rect 200264 79648 200942 79676
rect 200264 79636 200270 79648
rect 205634 79636 205640 79688
rect 205692 79676 205698 79688
rect 206434 79676 206462 79840
rect 224972 79824 225000 79852
rect 225368 79840 225374 79852
rect 225426 79840 225432 79892
rect 229784 79880 229790 79892
rect 229112 79852 229790 79880
rect 229112 79824 229140 79852
rect 229784 79840 229790 79852
rect 229842 79840 229848 79892
rect 230888 79840 230894 79892
rect 230946 79840 230952 79892
rect 231256 79840 231262 79892
rect 231314 79840 231320 79892
rect 231854 79840 231860 79892
rect 231912 79880 231918 79892
rect 232360 79880 232366 79892
rect 231912 79852 232366 79880
rect 231912 79840 231918 79852
rect 232360 79840 232366 79852
rect 232418 79840 232424 79892
rect 232728 79840 232734 79892
rect 232786 79840 232792 79892
rect 238156 79880 238162 79892
rect 237392 79852 238162 79880
rect 208394 79772 208400 79824
rect 208452 79812 208458 79824
rect 208992 79812 208998 79824
rect 208452 79784 208998 79812
rect 208452 79772 208458 79784
rect 208992 79772 208998 79784
rect 209050 79772 209056 79824
rect 209774 79772 209780 79824
rect 209832 79812 209838 79824
rect 210832 79812 210838 79824
rect 209832 79784 210838 79812
rect 209832 79772 209838 79784
rect 210832 79772 210838 79784
rect 210890 79772 210896 79824
rect 213914 79772 213920 79824
rect 213972 79812 213978 79824
rect 215156 79812 215162 79824
rect 213972 79784 215162 79812
rect 213972 79772 213978 79784
rect 215156 79772 215162 79784
rect 215214 79772 215220 79824
rect 219434 79772 219440 79824
rect 219492 79812 219498 79824
rect 219940 79812 219946 79824
rect 219492 79784 219946 79812
rect 219492 79772 219498 79784
rect 219940 79772 219946 79784
rect 219998 79772 220004 79824
rect 220906 79772 220912 79824
rect 220964 79812 220970 79824
rect 221780 79812 221786 79824
rect 220964 79784 221786 79812
rect 220964 79772 220970 79784
rect 221780 79772 221786 79784
rect 221838 79772 221844 79824
rect 222286 79772 222292 79824
rect 222344 79812 222350 79824
rect 223252 79812 223258 79824
rect 222344 79784 223258 79812
rect 222344 79772 222350 79784
rect 223252 79772 223258 79784
rect 223310 79772 223316 79824
rect 224954 79772 224960 79824
rect 225012 79772 225018 79824
rect 225046 79772 225052 79824
rect 225104 79812 225110 79824
rect 226104 79812 226110 79824
rect 225104 79784 226110 79812
rect 225104 79772 225110 79784
rect 226104 79772 226110 79784
rect 226162 79772 226168 79824
rect 227714 79772 227720 79824
rect 227772 79812 227778 79824
rect 228680 79812 228686 79824
rect 227772 79784 228686 79812
rect 227772 79772 227778 79784
rect 228680 79772 228686 79784
rect 228738 79772 228744 79824
rect 229094 79772 229100 79824
rect 229152 79772 229158 79824
rect 230906 79744 230934 79840
rect 230492 79716 230934 79744
rect 230492 79688 230520 79716
rect 205692 79648 206462 79676
rect 205692 79636 205698 79648
rect 224862 79636 224868 79688
rect 224920 79676 224926 79688
rect 225230 79676 225236 79688
rect 224920 79648 225236 79676
rect 224920 79636 224926 79648
rect 225230 79636 225236 79648
rect 225288 79636 225294 79688
rect 230474 79636 230480 79688
rect 230532 79636 230538 79688
rect 230566 79636 230572 79688
rect 230624 79676 230630 79688
rect 231274 79676 231302 79840
rect 230624 79648 231302 79676
rect 230624 79636 230630 79648
rect 231946 79636 231952 79688
rect 232004 79676 232010 79688
rect 232746 79676 232774 79840
rect 237392 79688 237420 79852
rect 238156 79840 238162 79852
rect 238214 79840 238220 79892
rect 244274 79840 244280 79892
rect 244332 79880 244338 79892
rect 244780 79880 244786 79892
rect 244332 79852 244786 79880
rect 244332 79840 244338 79852
rect 244780 79840 244786 79852
rect 244838 79840 244844 79892
rect 248742 79840 248748 79892
rect 248800 79880 248806 79892
rect 249610 79880 249616 79892
rect 248800 79852 249616 79880
rect 248800 79840 248806 79852
rect 249610 79840 249616 79852
rect 249668 79840 249674 79892
rect 251174 79840 251180 79892
rect 251232 79880 251238 79892
rect 251680 79880 251686 79892
rect 251232 79852 251686 79880
rect 251232 79840 251238 79852
rect 251680 79840 251686 79852
rect 251738 79840 251744 79892
rect 252646 79840 252652 79892
rect 252704 79880 252710 79892
rect 253520 79880 253526 79892
rect 252704 79852 253526 79880
rect 252704 79840 252710 79852
rect 253520 79840 253526 79852
rect 253578 79840 253584 79892
rect 254118 79840 254124 79892
rect 254176 79880 254182 79892
rect 254992 79880 254998 79892
rect 254176 79852 254998 79880
rect 254176 79840 254182 79852
rect 254992 79840 254998 79852
rect 255050 79840 255056 79892
rect 238754 79772 238760 79824
rect 238812 79812 238818 79824
rect 239628 79812 239634 79824
rect 238812 79784 239634 79812
rect 238812 79772 238818 79784
rect 239628 79772 239634 79784
rect 239686 79772 239692 79824
rect 241698 79772 241704 79824
rect 241756 79812 241762 79824
rect 242572 79812 242578 79824
rect 241756 79784 242578 79812
rect 241756 79772 241762 79784
rect 242572 79772 242578 79784
rect 242630 79772 242636 79824
rect 248414 79772 248420 79824
rect 248472 79812 248478 79824
rect 249104 79812 249110 79824
rect 248472 79784 249110 79812
rect 248472 79772 248478 79784
rect 249104 79772 249110 79784
rect 249162 79772 249168 79824
rect 252554 79772 252560 79824
rect 252612 79812 252618 79824
rect 253152 79812 253158 79824
rect 252612 79784 253158 79812
rect 252612 79772 252618 79784
rect 253152 79772 253158 79784
rect 253210 79772 253216 79824
rect 254026 79772 254032 79824
rect 254084 79812 254090 79824
rect 254624 79812 254630 79824
rect 254084 79784 254630 79812
rect 254084 79772 254090 79784
rect 254624 79772 254630 79784
rect 254682 79772 254688 79824
rect 256786 79772 256792 79824
rect 256844 79812 256850 79824
rect 257936 79812 257942 79824
rect 256844 79784 257942 79812
rect 256844 79772 256850 79784
rect 257936 79772 257942 79784
rect 257994 79772 258000 79824
rect 258074 79772 258080 79824
rect 258132 79812 258138 79824
rect 258672 79812 258678 79824
rect 258132 79784 258678 79812
rect 258132 79772 258138 79784
rect 258672 79772 258678 79784
rect 258730 79772 258736 79824
rect 232004 79648 232774 79676
rect 232004 79636 232010 79648
rect 237374 79636 237380 79688
rect 237432 79636 237438 79688
rect 80330 78752 80336 78804
rect 80388 78792 80394 78804
rect 447778 78792 447784 78804
rect 80388 78764 447784 78792
rect 80388 78752 80394 78764
rect 447778 78752 447784 78764
rect 447836 78752 447842 78804
rect 80238 78684 80244 78736
rect 80296 78724 80302 78736
rect 447870 78724 447876 78736
rect 80296 78696 447876 78724
rect 80296 78684 80302 78696
rect 447870 78684 447876 78696
rect 447928 78684 447934 78736
rect 112162 78616 112168 78668
rect 112220 78656 112226 78668
rect 114554 78656 114560 78668
rect 112220 78628 114560 78656
rect 112220 78616 112226 78628
rect 114554 78616 114560 78628
rect 114612 78616 114618 78668
rect 189626 78616 189632 78668
rect 189684 78656 189690 78668
rect 191374 78656 191380 78668
rect 189684 78628 191380 78656
rect 189684 78616 189690 78628
rect 191374 78616 191380 78628
rect 191432 78616 191438 78668
rect 97258 78548 97264 78600
rect 97316 78588 97322 78600
rect 105262 78588 105268 78600
rect 97316 78560 105268 78588
rect 97316 78548 97322 78560
rect 105262 78548 105268 78560
rect 105320 78548 105326 78600
rect 188522 78548 188528 78600
rect 188580 78588 188586 78600
rect 192570 78588 192576 78600
rect 188580 78560 192576 78588
rect 188580 78548 188586 78560
rect 192570 78548 192576 78560
rect 192628 78548 192634 78600
rect 70394 78480 70400 78532
rect 70452 78520 70458 78532
rect 101950 78520 101956 78532
rect 70452 78492 101956 78520
rect 70452 78480 70458 78492
rect 101950 78480 101956 78492
rect 102008 78480 102014 78532
rect 131574 78480 131580 78532
rect 131632 78520 131638 78532
rect 134518 78520 134524 78532
rect 131632 78492 134524 78520
rect 131632 78480 131638 78492
rect 134518 78480 134524 78492
rect 134576 78480 134582 78532
rect 185670 78480 185676 78532
rect 185728 78520 185734 78532
rect 191282 78520 191288 78532
rect 185728 78492 191288 78520
rect 185728 78480 185734 78492
rect 191282 78480 191288 78492
rect 191340 78480 191346 78532
rect 204990 78480 204996 78532
rect 205048 78520 205054 78532
rect 210418 78520 210424 78532
rect 205048 78492 210424 78520
rect 205048 78480 205054 78492
rect 210418 78480 210424 78492
rect 210476 78480 210482 78532
rect 65518 78412 65524 78464
rect 65576 78452 65582 78464
rect 99742 78452 99748 78464
rect 65576 78424 99748 78452
rect 65576 78412 65582 78424
rect 99742 78412 99748 78424
rect 99800 78412 99806 78464
rect 53098 78344 53104 78396
rect 53156 78384 53162 78396
rect 93210 78384 93216 78396
rect 53156 78356 93216 78384
rect 53156 78344 53162 78356
rect 93210 78344 93216 78356
rect 93268 78344 93274 78396
rect 110414 78344 110420 78396
rect 110472 78384 110478 78396
rect 114002 78384 114008 78396
rect 110472 78356 114008 78384
rect 110472 78344 110478 78356
rect 114002 78344 114008 78356
rect 114060 78344 114066 78396
rect 50338 78276 50344 78328
rect 50396 78316 50402 78328
rect 91094 78316 91100 78328
rect 50396 78288 91100 78316
rect 50396 78276 50402 78288
rect 91094 78276 91100 78288
rect 91152 78276 91158 78328
rect 93118 78276 93124 78328
rect 93176 78316 93182 78328
rect 96430 78316 96436 78328
rect 93176 78288 96436 78316
rect 93176 78276 93182 78288
rect 96430 78276 96436 78288
rect 96488 78276 96494 78328
rect 227990 78276 227996 78328
rect 228048 78316 228054 78328
rect 258718 78316 258724 78328
rect 228048 78288 258724 78316
rect 228048 78276 228054 78288
rect 258718 78276 258724 78288
rect 258776 78276 258782 78328
rect 28258 78208 28264 78260
rect 28316 78248 28322 78260
rect 86218 78248 86224 78260
rect 28316 78220 86224 78248
rect 28316 78208 28322 78220
rect 86218 78208 86224 78220
rect 86276 78208 86282 78260
rect 110506 78208 110512 78260
rect 110564 78248 110570 78260
rect 111058 78248 111064 78260
rect 110564 78220 111064 78248
rect 110564 78208 110570 78220
rect 111058 78208 111064 78220
rect 111116 78208 111122 78260
rect 207198 78208 207204 78260
rect 207256 78248 207262 78260
rect 213086 78248 213092 78260
rect 207256 78220 213092 78248
rect 207256 78208 207262 78220
rect 213086 78208 213092 78220
rect 213144 78208 213150 78260
rect 226886 78208 226892 78260
rect 226944 78248 226950 78260
rect 289078 78248 289084 78260
rect 226944 78220 289084 78248
rect 226944 78208 226950 78220
rect 289078 78208 289084 78220
rect 289136 78208 289142 78260
rect 32398 78140 32404 78192
rect 32456 78180 32462 78192
rect 88794 78180 88800 78192
rect 32456 78152 88800 78180
rect 32456 78140 32462 78152
rect 88794 78140 88800 78152
rect 88852 78140 88858 78192
rect 136358 78140 136364 78192
rect 136416 78180 136422 78192
rect 166442 78180 166448 78192
rect 136416 78152 166448 78180
rect 136416 78140 136422 78152
rect 166442 78140 166448 78152
rect 166500 78140 166506 78192
rect 215938 78140 215944 78192
rect 215996 78180 216002 78192
rect 226978 78180 226984 78192
rect 215996 78152 226984 78180
rect 215996 78140 216002 78152
rect 226978 78140 226984 78152
rect 227036 78140 227042 78192
rect 259086 78140 259092 78192
rect 259144 78180 259150 78192
rect 418798 78180 418804 78192
rect 259144 78152 418804 78180
rect 259144 78140 259150 78152
rect 418798 78140 418804 78152
rect 418856 78140 418862 78192
rect 25498 78072 25504 78124
rect 25556 78112 25562 78124
rect 85942 78112 85948 78124
rect 25556 78084 85948 78112
rect 25556 78072 25562 78084
rect 85942 78072 85948 78084
rect 86000 78072 86006 78124
rect 101398 78072 101404 78124
rect 101456 78112 101462 78124
rect 106274 78112 106280 78124
rect 101456 78084 106280 78112
rect 101456 78072 101462 78084
rect 106274 78072 106280 78084
rect 106332 78072 106338 78124
rect 111058 78072 111064 78124
rect 111116 78112 111122 78124
rect 113634 78112 113640 78124
rect 111116 78084 113640 78112
rect 111116 78072 111122 78084
rect 113634 78072 113640 78084
rect 113692 78072 113698 78124
rect 129366 78072 129372 78124
rect 129424 78112 129430 78124
rect 135898 78112 135904 78124
rect 129424 78084 135904 78112
rect 129424 78072 129430 78084
rect 135898 78072 135904 78084
rect 135956 78072 135962 78124
rect 153838 78072 153844 78124
rect 153896 78112 153902 78124
rect 188338 78112 188344 78124
rect 153896 78084 188344 78112
rect 153896 78072 153902 78084
rect 188338 78072 188344 78084
rect 188396 78072 188402 78124
rect 209406 78072 209412 78124
rect 209464 78112 209470 78124
rect 214558 78112 214564 78124
rect 209464 78084 214564 78112
rect 209464 78072 209470 78084
rect 214558 78072 214564 78084
rect 214616 78072 214622 78124
rect 220354 78072 220360 78124
rect 220412 78112 220418 78124
rect 255958 78112 255964 78124
rect 220412 78084 255964 78112
rect 220412 78072 220418 78084
rect 255958 78072 255964 78084
rect 256016 78072 256022 78124
rect 260098 78072 260104 78124
rect 260156 78112 260162 78124
rect 422938 78112 422944 78124
rect 260156 78084 422944 78112
rect 260156 78072 260162 78084
rect 422938 78072 422944 78084
rect 422996 78072 423002 78124
rect 15838 78004 15844 78056
rect 15896 78044 15902 78056
rect 83274 78044 83280 78056
rect 15896 78016 83280 78044
rect 15896 78004 15902 78016
rect 83274 78004 83280 78016
rect 83332 78004 83338 78056
rect 120626 78004 120632 78056
rect 120684 78044 120690 78056
rect 126238 78044 126244 78056
rect 120684 78016 126244 78044
rect 120684 78004 120690 78016
rect 126238 78004 126244 78016
rect 126296 78004 126302 78056
rect 149514 78004 149520 78056
rect 149572 78044 149578 78056
rect 187050 78044 187056 78056
rect 149572 78016 187056 78044
rect 149572 78004 149578 78016
rect 187050 78004 187056 78016
rect 187108 78004 187114 78056
rect 198458 78004 198464 78056
rect 198516 78044 198522 78056
rect 203518 78044 203524 78056
rect 198516 78016 203524 78044
rect 198516 78004 198522 78016
rect 203518 78004 203524 78016
rect 203576 78004 203582 78056
rect 208302 78004 208308 78056
rect 208360 78044 208366 78056
rect 213178 78044 213184 78056
rect 208360 78016 213184 78044
rect 208360 78004 208366 78016
rect 213178 78004 213184 78016
rect 213236 78004 213242 78056
rect 222562 78004 222568 78056
rect 222620 78044 222626 78056
rect 407758 78044 407764 78056
rect 222620 78016 407764 78044
rect 222620 78004 222626 78016
rect 407758 78004 407764 78016
rect 407816 78004 407822 78056
rect 10318 77936 10324 77988
rect 10376 77976 10382 77988
rect 81434 77976 81440 77988
rect 10376 77948 81440 77976
rect 10376 77936 10382 77948
rect 81434 77936 81440 77948
rect 81492 77936 81498 77988
rect 102134 77936 102140 77988
rect 102192 77976 102198 77988
rect 111794 77976 111800 77988
rect 102192 77948 111800 77976
rect 102192 77936 102198 77948
rect 111794 77936 111800 77948
rect 111852 77936 111858 77988
rect 131942 77936 131948 77988
rect 132000 77976 132006 77988
rect 141418 77976 141424 77988
rect 132000 77948 141424 77976
rect 132000 77936 132006 77948
rect 141418 77936 141424 77948
rect 141476 77936 141482 77988
rect 143994 77936 144000 77988
rect 144052 77976 144058 77988
rect 186958 77976 186964 77988
rect 144052 77948 186964 77976
rect 144052 77936 144058 77948
rect 186958 77936 186964 77948
rect 187016 77936 187022 77988
rect 224678 77936 224684 77988
rect 224736 77976 224742 77988
rect 411898 77976 411904 77988
rect 224736 77948 411904 77976
rect 224736 77936 224742 77948
rect 411898 77936 411904 77948
rect 411956 77936 411962 77988
rect 124214 77868 124220 77920
rect 124272 77908 124278 77920
rect 129090 77908 129096 77920
rect 124272 77880 129096 77908
rect 124272 77868 124278 77880
rect 129090 77868 129096 77880
rect 129148 77868 129154 77920
rect 107654 77800 107660 77852
rect 107712 77840 107718 77852
rect 113266 77840 113272 77852
rect 107712 77812 113272 77840
rect 107712 77800 107718 77812
rect 113266 77800 113272 77812
rect 113324 77800 113330 77852
rect 121362 77800 121368 77852
rect 121420 77840 121426 77852
rect 123478 77840 123484 77852
rect 121420 77812 123484 77840
rect 121420 77800 121426 77812
rect 123478 77800 123484 77812
rect 123536 77800 123542 77852
rect 118418 77732 118424 77784
rect 118476 77772 118482 77784
rect 124214 77772 124220 77784
rect 118476 77744 124220 77772
rect 118476 77732 118482 77744
rect 124214 77732 124220 77744
rect 124272 77732 124278 77784
rect 190730 77664 190736 77716
rect 190788 77704 190794 77716
rect 192386 77704 192392 77716
rect 190788 77676 192392 77704
rect 190788 77664 190794 77676
rect 192386 77664 192392 77676
rect 192444 77664 192450 77716
rect 106918 77460 106924 77512
rect 106976 77500 106982 77512
rect 108850 77500 108856 77512
rect 106976 77472 108856 77500
rect 106976 77460 106982 77472
rect 108850 77460 108856 77472
rect 108908 77460 108914 77512
rect 144178 77500 144184 77512
rect 142126 77472 144184 77500
rect 105538 77392 105544 77444
rect 105596 77432 105602 77444
rect 107378 77432 107384 77444
rect 105596 77404 107384 77432
rect 105596 77392 105602 77404
rect 107378 77392 107384 77404
rect 107436 77392 107442 77444
rect 135622 77392 135628 77444
rect 135680 77432 135686 77444
rect 142126 77432 142154 77472
rect 144178 77460 144184 77472
rect 144236 77460 144242 77512
rect 201678 77460 201684 77512
rect 201736 77500 201742 77512
rect 209038 77500 209044 77512
rect 201736 77472 209044 77500
rect 201736 77460 201742 77472
rect 209038 77460 209044 77472
rect 209096 77460 209102 77512
rect 135680 77404 142154 77432
rect 135680 77392 135686 77404
rect 142430 77392 142436 77444
rect 142488 77392 142494 77444
rect 187510 77392 187516 77444
rect 187568 77432 187574 77444
rect 191098 77432 191104 77444
rect 187568 77404 191104 77432
rect 187568 77392 187574 77404
rect 191098 77392 191104 77404
rect 191156 77392 191162 77444
rect 202782 77392 202788 77444
rect 202840 77432 202846 77444
rect 207750 77432 207756 77444
rect 202840 77404 207756 77432
rect 202840 77392 202846 77404
rect 207750 77392 207756 77404
rect 207808 77392 207814 77444
rect 229186 77392 229192 77444
rect 229244 77392 229250 77444
rect 100018 77324 100024 77376
rect 100076 77364 100082 77376
rect 103054 77364 103060 77376
rect 100076 77336 103060 77364
rect 100076 77324 100082 77336
rect 103054 77324 103060 77336
rect 103112 77324 103118 77376
rect 107010 77324 107016 77376
rect 107068 77364 107074 77376
rect 108482 77364 108488 77376
rect 107068 77336 108488 77364
rect 107068 77324 107074 77336
rect 108482 77324 108488 77336
rect 108540 77324 108546 77376
rect 118050 77324 118056 77376
rect 118108 77364 118114 77376
rect 119338 77364 119344 77376
rect 118108 77336 119344 77364
rect 118108 77324 118114 77336
rect 119338 77324 119344 77336
rect 119396 77324 119402 77376
rect 123202 77324 123208 77376
rect 123260 77364 123266 77376
rect 128998 77364 129004 77376
rect 123260 77336 129004 77364
rect 123260 77324 123266 77336
rect 128998 77324 129004 77336
rect 129056 77324 129062 77376
rect 135346 77324 135352 77376
rect 135404 77364 135410 77376
rect 137278 77364 137284 77376
rect 135404 77336 137284 77364
rect 135404 77324 135410 77336
rect 137278 77324 137284 77336
rect 137336 77324 137342 77376
rect 81526 77256 81532 77308
rect 81584 77296 81590 77308
rect 82538 77296 82544 77308
rect 81584 77268 82544 77296
rect 81584 77256 81590 77268
rect 82538 77256 82544 77268
rect 82596 77256 82602 77308
rect 82906 77256 82912 77308
rect 82964 77296 82970 77308
rect 84010 77296 84016 77308
rect 82964 77268 84016 77296
rect 82964 77256 82970 77268
rect 84010 77256 84016 77268
rect 84068 77256 84074 77308
rect 86954 77256 86960 77308
rect 87012 77296 87018 77308
rect 87230 77296 87236 77308
rect 87012 77268 87236 77296
rect 87012 77256 87018 77268
rect 87230 77256 87236 77268
rect 87288 77256 87294 77308
rect 88518 77256 88524 77308
rect 88576 77296 88582 77308
rect 89530 77296 89536 77308
rect 88576 77268 89536 77296
rect 88576 77256 88582 77268
rect 89530 77256 89536 77268
rect 89588 77256 89594 77308
rect 93946 77256 93952 77308
rect 94004 77296 94010 77308
rect 94130 77296 94136 77308
rect 94004 77268 94136 77296
rect 94004 77256 94010 77268
rect 94130 77256 94136 77268
rect 94188 77256 94194 77308
rect 100846 77256 100852 77308
rect 100904 77296 100910 77308
rect 101582 77296 101588 77308
rect 100904 77268 101588 77296
rect 100904 77256 100910 77268
rect 101582 77256 101588 77268
rect 101640 77256 101646 77308
rect 104986 77256 104992 77308
rect 105044 77296 105050 77308
rect 105906 77296 105912 77308
rect 105044 77268 105912 77296
rect 105044 77256 105050 77268
rect 105906 77256 105912 77268
rect 105964 77256 105970 77308
rect 107746 77256 107752 77308
rect 107804 77296 107810 77308
rect 108114 77296 108120 77308
rect 107804 77268 108120 77296
rect 107804 77256 107810 77268
rect 108114 77256 108120 77268
rect 108172 77256 108178 77308
rect 108298 77256 108304 77308
rect 108356 77296 108362 77308
rect 109586 77296 109592 77308
rect 108356 77268 109592 77296
rect 108356 77256 108362 77268
rect 109586 77256 109592 77268
rect 109644 77256 109650 77308
rect 109678 77256 109684 77308
rect 109736 77296 109742 77308
rect 110690 77296 110696 77308
rect 109736 77268 110696 77296
rect 109736 77256 109742 77268
rect 110690 77256 110696 77268
rect 110748 77256 110754 77308
rect 111886 77256 111892 77308
rect 111944 77296 111950 77308
rect 112898 77296 112904 77308
rect 111944 77268 112904 77296
rect 111944 77256 111950 77268
rect 112898 77256 112904 77268
rect 112956 77256 112962 77308
rect 118786 77256 118792 77308
rect 118844 77296 118850 77308
rect 119798 77296 119804 77308
rect 118844 77268 119804 77296
rect 118844 77256 118850 77268
rect 119798 77256 119804 77268
rect 119856 77256 119862 77308
rect 120994 77256 121000 77308
rect 121052 77296 121058 77308
rect 122098 77296 122104 77308
rect 121052 77268 122104 77296
rect 121052 77256 121058 77268
rect 122098 77256 122104 77268
rect 122156 77256 122162 77308
rect 125778 77256 125784 77308
rect 125836 77296 125842 77308
rect 126422 77296 126428 77308
rect 125836 77268 126428 77296
rect 125836 77256 125842 77268
rect 126422 77256 126428 77268
rect 126480 77256 126486 77308
rect 127986 77256 127992 77308
rect 128044 77296 128050 77308
rect 129182 77296 129188 77308
rect 128044 77268 129188 77296
rect 128044 77256 128050 77268
rect 129182 77256 129188 77268
rect 129240 77256 129246 77308
rect 129734 77256 129740 77308
rect 129792 77296 129798 77308
rect 130378 77296 130384 77308
rect 129792 77268 130384 77296
rect 129792 77256 129798 77268
rect 130378 77256 130384 77268
rect 130436 77256 130442 77308
rect 132678 77256 132684 77308
rect 132736 77296 132742 77308
rect 133322 77296 133328 77308
rect 132736 77268 133328 77296
rect 132736 77256 132742 77268
rect 133322 77256 133328 77268
rect 133380 77256 133386 77308
rect 136726 77256 136732 77308
rect 136784 77296 136790 77308
rect 137370 77296 137376 77308
rect 136784 77268 137376 77296
rect 136784 77256 136790 77268
rect 137370 77256 137376 77268
rect 137428 77256 137434 77308
rect 138198 77256 138204 77308
rect 138256 77296 138262 77308
rect 139210 77296 139216 77308
rect 138256 77268 139216 77296
rect 138256 77256 138262 77268
rect 139210 77256 139216 77268
rect 139268 77256 139274 77308
rect 139486 77256 139492 77308
rect 139544 77296 139550 77308
rect 140590 77296 140596 77308
rect 139544 77268 140596 77296
rect 139544 77256 139550 77268
rect 140590 77256 140596 77268
rect 140648 77256 140654 77308
rect 93854 77188 93860 77240
rect 93912 77228 93918 77240
rect 94958 77228 94964 77240
rect 93912 77200 94964 77228
rect 93912 77188 93918 77200
rect 94958 77188 94964 77200
rect 95016 77188 95022 77240
rect 109218 77188 109224 77240
rect 109276 77228 109282 77240
rect 109954 77228 109960 77240
rect 109276 77200 109960 77228
rect 109276 77188 109282 77200
rect 109954 77188 109960 77200
rect 110012 77188 110018 77240
rect 125686 77188 125692 77240
rect 125744 77228 125750 77240
rect 126790 77228 126796 77240
rect 125744 77200 126796 77228
rect 125744 77188 125750 77200
rect 126790 77188 126796 77200
rect 126848 77188 126854 77240
rect 132586 77188 132592 77240
rect 132644 77228 132650 77240
rect 133690 77228 133696 77240
rect 132644 77200 133696 77228
rect 132644 77188 132650 77200
rect 133690 77188 133696 77200
rect 133748 77188 133754 77240
rect 136634 77188 136640 77240
rect 136692 77228 136698 77240
rect 137738 77228 137744 77240
rect 136692 77200 137744 77228
rect 136692 77188 136698 77200
rect 137738 77188 137744 77200
rect 137796 77188 137802 77240
rect 138106 77188 138112 77240
rect 138164 77228 138170 77240
rect 138842 77228 138848 77240
rect 138164 77200 138848 77228
rect 138164 77188 138170 77200
rect 138842 77188 138848 77200
rect 138900 77188 138906 77240
rect 87138 77120 87144 77172
rect 87196 77160 87202 77172
rect 87690 77160 87696 77172
rect 87196 77132 87696 77160
rect 87196 77120 87202 77132
rect 87690 77120 87696 77132
rect 87748 77120 87754 77172
rect 92566 77120 92572 77172
rect 92624 77160 92630 77172
rect 93486 77160 93492 77172
rect 92624 77132 93492 77160
rect 92624 77120 92630 77132
rect 93486 77120 93492 77132
rect 93544 77120 93550 77172
rect 93946 77120 93952 77172
rect 94004 77160 94010 77172
rect 94590 77160 94596 77172
rect 94004 77132 94596 77160
rect 94004 77120 94010 77132
rect 94590 77120 94596 77132
rect 94648 77120 94654 77172
rect 110690 77120 110696 77172
rect 110748 77160 110754 77172
rect 111426 77160 111432 77172
rect 110748 77132 111432 77160
rect 110748 77120 110754 77132
rect 111426 77120 111432 77132
rect 111484 77120 111490 77172
rect 142448 77104 142476 77392
rect 167178 77324 167184 77376
rect 167236 77364 167242 77376
rect 169018 77364 169024 77376
rect 167236 77336 169024 77364
rect 167236 77324 167242 77336
rect 169018 77324 169024 77336
rect 169076 77324 169082 77376
rect 192938 77324 192944 77376
rect 192996 77364 193002 77376
rect 193858 77364 193864 77376
rect 192996 77336 193864 77364
rect 192996 77324 193002 77336
rect 193858 77324 193864 77336
rect 193916 77324 193922 77376
rect 194042 77324 194048 77376
rect 194100 77364 194106 77376
rect 195238 77364 195244 77376
rect 194100 77336 195244 77364
rect 194100 77324 194106 77336
rect 195238 77324 195244 77336
rect 195296 77324 195302 77376
rect 206094 77324 206100 77376
rect 206152 77364 206158 77376
rect 209130 77364 209136 77376
rect 206152 77336 209136 77364
rect 206152 77324 206158 77336
rect 209130 77324 209136 77336
rect 209188 77324 209194 77376
rect 210510 77324 210516 77376
rect 210568 77364 210574 77376
rect 217318 77364 217324 77376
rect 210568 77336 217324 77364
rect 210568 77324 210574 77336
rect 217318 77324 217324 77336
rect 217376 77324 217382 77376
rect 143626 77256 143632 77308
rect 143684 77296 143690 77308
rect 144638 77296 144644 77308
rect 143684 77268 144644 77296
rect 143684 77256 143690 77268
rect 144638 77256 144644 77268
rect 144696 77256 144702 77308
rect 145098 77256 145104 77308
rect 145156 77296 145162 77308
rect 145742 77296 145748 77308
rect 145156 77268 145748 77296
rect 145156 77256 145162 77268
rect 145742 77256 145748 77268
rect 145800 77256 145806 77308
rect 147674 77256 147680 77308
rect 147732 77296 147738 77308
rect 148318 77296 148324 77308
rect 147732 77268 148324 77296
rect 147732 77256 147738 77268
rect 148318 77256 148324 77268
rect 148376 77256 148382 77308
rect 149054 77256 149060 77308
rect 149112 77296 149118 77308
rect 150158 77296 150164 77308
rect 149112 77268 150164 77296
rect 149112 77256 149118 77268
rect 150158 77256 150164 77268
rect 150216 77256 150222 77308
rect 150618 77256 150624 77308
rect 150676 77296 150682 77308
rect 151630 77296 151636 77308
rect 150676 77268 151636 77296
rect 150676 77256 150682 77268
rect 151630 77256 151636 77268
rect 151688 77256 151694 77308
rect 154574 77256 154580 77308
rect 154632 77296 154638 77308
rect 155586 77296 155592 77308
rect 154632 77268 155592 77296
rect 154632 77256 154638 77268
rect 155586 77256 155592 77268
rect 155644 77256 155650 77308
rect 155954 77256 155960 77308
rect 156012 77296 156018 77308
rect 156690 77296 156696 77308
rect 156012 77268 156696 77296
rect 156012 77256 156018 77268
rect 156690 77256 156696 77268
rect 156748 77256 156754 77308
rect 168466 77256 168472 77308
rect 168524 77296 168530 77308
rect 169478 77296 169484 77308
rect 168524 77268 169484 77296
rect 168524 77256 168530 77268
rect 169478 77256 169484 77268
rect 169536 77256 169542 77308
rect 175366 77256 175372 77308
rect 175424 77296 175430 77308
rect 176378 77296 176384 77308
rect 175424 77268 176384 77296
rect 175424 77256 175430 77268
rect 176378 77256 176384 77268
rect 176436 77256 176442 77308
rect 191834 77256 191840 77308
rect 191892 77296 191898 77308
rect 192018 77296 192024 77308
rect 191892 77268 192024 77296
rect 191892 77256 191898 77268
rect 192018 77256 192024 77268
rect 192076 77256 192082 77308
rect 193214 77256 193220 77308
rect 193272 77296 193278 77308
rect 193582 77296 193588 77308
rect 193272 77268 193588 77296
rect 193272 77256 193278 77268
rect 193582 77256 193588 77268
rect 193640 77256 193646 77308
rect 194686 77256 194692 77308
rect 194744 77296 194750 77308
rect 195054 77296 195060 77308
rect 194744 77268 195060 77296
rect 194744 77256 194750 77268
rect 195054 77256 195060 77268
rect 195112 77256 195118 77308
rect 198734 77256 198740 77308
rect 198792 77296 198798 77308
rect 199470 77296 199476 77308
rect 198792 77268 199476 77296
rect 198792 77256 198798 77268
rect 199470 77256 199476 77268
rect 199528 77256 199534 77308
rect 203886 77256 203892 77308
rect 203944 77296 203950 77308
rect 206278 77296 206284 77308
rect 203944 77268 206284 77296
rect 203944 77256 203950 77268
rect 206278 77256 206284 77268
rect 206336 77256 206342 77308
rect 211246 77256 211252 77308
rect 211304 77296 211310 77308
rect 211522 77296 211528 77308
rect 211304 77268 211528 77296
rect 211304 77256 211310 77268
rect 211522 77256 211528 77268
rect 211580 77256 211586 77308
rect 212626 77256 212632 77308
rect 212684 77296 212690 77308
rect 213270 77296 213276 77308
rect 212684 77268 213276 77296
rect 212684 77256 212690 77268
rect 213270 77256 213276 77268
rect 213328 77256 213334 77308
rect 213730 77256 213736 77308
rect 213788 77296 213794 77308
rect 215938 77296 215944 77308
rect 213788 77268 215944 77296
rect 213788 77256 213794 77268
rect 215938 77256 215944 77268
rect 215996 77256 216002 77308
rect 218146 77256 218152 77308
rect 218204 77296 218210 77308
rect 218330 77296 218336 77308
rect 218204 77268 218336 77296
rect 218204 77256 218210 77268
rect 218330 77256 218336 77268
rect 218388 77256 218394 77308
rect 219526 77256 219532 77308
rect 219584 77296 219590 77308
rect 220630 77296 220636 77308
rect 219584 77268 220636 77296
rect 219584 77256 219590 77268
rect 220630 77256 220636 77268
rect 220688 77256 220694 77308
rect 223666 77256 223672 77308
rect 223724 77296 223730 77308
rect 223850 77296 223856 77308
rect 223724 77268 223856 77296
rect 223724 77256 223730 77268
rect 223850 77256 223856 77268
rect 223908 77256 223914 77308
rect 226426 77256 226432 77308
rect 226484 77296 226490 77308
rect 227530 77296 227536 77308
rect 226484 77268 227536 77296
rect 226484 77256 226490 77268
rect 227530 77256 227536 77268
rect 227588 77256 227594 77308
rect 150526 77188 150532 77240
rect 150584 77228 150590 77240
rect 151262 77228 151268 77240
rect 150584 77200 151268 77228
rect 150584 77188 150590 77200
rect 151262 77188 151268 77200
rect 151320 77188 151326 77240
rect 168374 77188 168380 77240
rect 168432 77228 168438 77240
rect 169110 77228 169116 77240
rect 168432 77200 169116 77228
rect 168432 77188 168438 77200
rect 169110 77188 169116 77200
rect 169168 77188 169174 77240
rect 211154 77188 211160 77240
rect 211212 77228 211218 77240
rect 211706 77228 211712 77240
rect 211212 77200 211712 77228
rect 211212 77188 211218 77200
rect 211706 77188 211712 77200
rect 211764 77188 211770 77240
rect 214098 77188 214104 77240
rect 214156 77228 214162 77240
rect 214742 77228 214748 77240
rect 214156 77200 214748 77228
rect 214156 77188 214162 77200
rect 214742 77188 214748 77200
rect 214800 77188 214806 77240
rect 218054 77188 218060 77240
rect 218112 77228 218118 77240
rect 219158 77228 219164 77240
rect 218112 77200 219164 77228
rect 218112 77188 218118 77200
rect 219158 77188 219164 77200
rect 219216 77188 219222 77240
rect 223574 77188 223580 77240
rect 223632 77228 223638 77240
rect 224218 77228 224224 77240
rect 223632 77200 224224 77228
rect 223632 77188 223638 77200
rect 224218 77188 224224 77200
rect 224276 77188 224282 77240
rect 226518 77188 226524 77240
rect 226576 77228 226582 77240
rect 227162 77228 227168 77240
rect 226576 77200 227168 77228
rect 226576 77188 226582 77200
rect 227162 77188 227168 77200
rect 227220 77188 227226 77240
rect 229204 77228 229232 77392
rect 242986 77324 242992 77376
rect 243044 77364 243050 77376
rect 243998 77364 244004 77376
rect 243044 77336 244004 77364
rect 243044 77324 243050 77336
rect 243998 77324 244004 77336
rect 244056 77324 244062 77376
rect 234614 77256 234620 77308
rect 234672 77296 234678 77308
rect 235626 77296 235632 77308
rect 234672 77268 235632 77296
rect 234672 77256 234678 77268
rect 235626 77256 235632 77268
rect 235684 77256 235690 77308
rect 236086 77256 236092 77308
rect 236144 77296 236150 77308
rect 236638 77296 236644 77308
rect 236144 77268 236644 77296
rect 236144 77256 236150 77268
rect 236638 77256 236644 77268
rect 236696 77256 236702 77308
rect 238938 77256 238944 77308
rect 238996 77296 239002 77308
rect 239950 77296 239956 77308
rect 238996 77268 239956 77296
rect 238996 77256 239002 77268
rect 239950 77256 239956 77268
rect 240008 77256 240014 77308
rect 240226 77256 240232 77308
rect 240284 77296 240290 77308
rect 241054 77296 241060 77308
rect 240284 77268 241060 77296
rect 240284 77256 240290 77268
rect 241054 77256 241060 77268
rect 241112 77256 241118 77308
rect 241514 77256 241520 77308
rect 241572 77296 241578 77308
rect 242158 77296 242164 77308
rect 241572 77268 242164 77296
rect 241572 77256 241578 77268
rect 242158 77256 242164 77268
rect 242216 77256 242222 77308
rect 243078 77256 243084 77308
rect 243136 77296 243142 77308
rect 243630 77296 243636 77308
rect 243136 77268 243636 77296
rect 243136 77256 243142 77268
rect 243630 77256 243636 77268
rect 243688 77256 243694 77308
rect 244458 77256 244464 77308
rect 244516 77296 244522 77308
rect 245470 77296 245476 77308
rect 244516 77268 245476 77296
rect 244516 77256 244522 77268
rect 245470 77256 245476 77268
rect 245528 77256 245534 77308
rect 245746 77256 245752 77308
rect 245804 77296 245810 77308
rect 246574 77296 246580 77308
rect 245804 77268 246580 77296
rect 245804 77256 245810 77268
rect 246574 77256 246580 77268
rect 246632 77256 246638 77308
rect 247126 77256 247132 77308
rect 247184 77296 247190 77308
rect 247678 77296 247684 77308
rect 247184 77268 247684 77296
rect 247184 77256 247190 77268
rect 247678 77256 247684 77268
rect 247736 77256 247742 77308
rect 248506 77256 248512 77308
rect 248564 77296 248570 77308
rect 249426 77296 249432 77308
rect 248564 77268 249432 77296
rect 248564 77256 248570 77268
rect 249426 77256 249432 77268
rect 249484 77256 249490 77308
rect 249794 77256 249800 77308
rect 249852 77296 249858 77308
rect 250346 77296 250352 77308
rect 249852 77268 250352 77296
rect 249852 77256 249858 77268
rect 250346 77256 250352 77268
rect 250404 77256 250410 77308
rect 251358 77256 251364 77308
rect 251416 77296 251422 77308
rect 252370 77296 252376 77308
rect 251416 77268 252376 77296
rect 251416 77256 251422 77268
rect 252370 77256 252376 77268
rect 252428 77256 252434 77308
rect 229278 77228 229284 77240
rect 229204 77200 229284 77228
rect 229278 77188 229284 77200
rect 229336 77188 229342 77240
rect 235994 77188 236000 77240
rect 236052 77228 236058 77240
rect 237006 77228 237012 77240
rect 236052 77200 237012 77228
rect 236052 77188 236058 77200
rect 237006 77188 237012 77200
rect 237064 77188 237070 77240
rect 242894 77188 242900 77240
rect 242952 77228 242958 77240
rect 243262 77228 243268 77240
rect 242952 77200 243268 77228
rect 242952 77188 242958 77200
rect 243262 77188 243268 77200
rect 243320 77188 243326 77240
rect 247034 77188 247040 77240
rect 247092 77228 247098 77240
rect 248046 77228 248052 77240
rect 247092 77200 248052 77228
rect 247092 77188 247098 77200
rect 248046 77188 248052 77200
rect 248104 77188 248110 77240
rect 191834 77120 191840 77172
rect 191892 77160 191898 77172
rect 192478 77160 192484 77172
rect 191892 77132 192484 77160
rect 191892 77120 191898 77132
rect 192478 77120 192484 77132
rect 192536 77120 192542 77172
rect 218146 77120 218152 77172
rect 218204 77160 218210 77172
rect 218790 77160 218796 77172
rect 218204 77132 218796 77160
rect 218204 77120 218210 77132
rect 218790 77120 218796 77132
rect 218848 77120 218854 77172
rect 142430 77052 142436 77104
rect 142488 77052 142494 77104
rect 255590 77052 255596 77104
rect 255648 77092 255654 77104
rect 256418 77092 256424 77104
rect 255648 77064 256424 77092
rect 255648 77052 255654 77064
rect 256418 77052 256424 77064
rect 256476 77052 256482 77104
rect 170030 76780 170036 76832
rect 170088 76820 170094 76832
rect 291194 76820 291200 76832
rect 170088 76792 291200 76820
rect 170088 76780 170094 76792
rect 291194 76780 291200 76792
rect 291252 76780 291258 76832
rect 216766 76712 216772 76764
rect 216824 76752 216830 76764
rect 441614 76752 441620 76764
rect 216824 76724 441620 76752
rect 216824 76712 216830 76724
rect 441614 76712 441620 76724
rect 441672 76712 441678 76764
rect 217778 76644 217784 76696
rect 217836 76684 217842 76696
rect 445754 76684 445760 76696
rect 217836 76656 445760 76684
rect 217836 76644 217842 76656
rect 445754 76644 445760 76656
rect 445812 76644 445818 76696
rect 51074 76576 51080 76628
rect 51132 76616 51138 76628
rect 95694 76616 95700 76628
rect 51132 76588 95700 76616
rect 51132 76576 51138 76588
rect 95694 76576 95700 76588
rect 95752 76576 95758 76628
rect 225230 76576 225236 76628
rect 225288 76616 225294 76628
rect 469214 76616 469220 76628
rect 225288 76588 469220 76616
rect 225288 76576 225294 76588
rect 469214 76576 469220 76588
rect 469272 76576 469278 76628
rect 49694 76508 49700 76560
rect 49752 76548 49758 76560
rect 95326 76548 95332 76560
rect 49752 76520 95332 76548
rect 49752 76508 49758 76520
rect 95326 76508 95332 76520
rect 95384 76508 95390 76560
rect 257614 76508 257620 76560
rect 257672 76548 257678 76560
rect 574094 76548 574100 76560
rect 257672 76520 574100 76548
rect 257672 76508 257678 76520
rect 574094 76508 574100 76520
rect 574152 76508 574158 76560
rect 86954 75624 86960 75676
rect 87012 75664 87018 75676
rect 88058 75664 88064 75676
rect 87012 75636 88064 75664
rect 87012 75624 87018 75636
rect 88058 75624 88064 75636
rect 88116 75624 88122 75676
rect 168834 75420 168840 75472
rect 168892 75460 168898 75472
rect 287054 75460 287060 75472
rect 168892 75432 287060 75460
rect 168892 75420 168898 75432
rect 287054 75420 287060 75432
rect 287112 75420 287118 75472
rect 195882 75352 195888 75404
rect 195940 75392 195946 75404
rect 373994 75392 374000 75404
rect 195940 75364 374000 75392
rect 195940 75352 195946 75364
rect 373994 75352 374000 75364
rect 374052 75352 374058 75404
rect 214466 75284 214472 75336
rect 214524 75324 214530 75336
rect 434714 75324 434720 75336
rect 214524 75296 434720 75324
rect 214524 75284 214530 75296
rect 434714 75284 434720 75296
rect 434772 75284 434778 75336
rect 215570 75216 215576 75268
rect 215628 75256 215634 75268
rect 438854 75256 438860 75268
rect 215628 75228 438860 75256
rect 215628 75216 215634 75228
rect 438854 75216 438860 75228
rect 438912 75216 438918 75268
rect 37274 75148 37280 75200
rect 37332 75188 37338 75200
rect 91738 75188 91744 75200
rect 37332 75160 91744 75188
rect 37332 75148 37338 75160
rect 91738 75148 91744 75160
rect 91796 75148 91802 75200
rect 161566 75148 161572 75200
rect 161624 75188 161630 75200
rect 162578 75188 162584 75200
rect 161624 75160 162584 75188
rect 161624 75148 161630 75160
rect 162578 75148 162584 75160
rect 162636 75148 162642 75200
rect 162946 75148 162952 75200
rect 163004 75188 163010 75200
rect 164050 75188 164056 75200
rect 163004 75160 164056 75188
rect 163004 75148 163010 75160
rect 164050 75148 164056 75160
rect 164108 75148 164114 75200
rect 164326 75148 164332 75200
rect 164384 75188 164390 75200
rect 165062 75188 165068 75200
rect 164384 75160 165068 75188
rect 164384 75148 164390 75160
rect 165062 75148 165068 75160
rect 165120 75148 165126 75200
rect 176838 75148 176844 75200
rect 176896 75188 176902 75200
rect 177850 75188 177856 75200
rect 176896 75160 177856 75188
rect 176896 75148 176902 75160
rect 177850 75148 177856 75160
rect 177908 75148 177914 75200
rect 180794 75148 180800 75200
rect 180852 75188 180858 75200
rect 181898 75188 181904 75200
rect 180852 75160 181904 75188
rect 180852 75148 180858 75160
rect 181898 75148 181904 75160
rect 181956 75148 181962 75200
rect 182358 75148 182364 75200
rect 182416 75188 182422 75200
rect 183370 75188 183376 75200
rect 182416 75160 183376 75188
rect 182416 75148 182422 75160
rect 183370 75148 183376 75160
rect 183428 75148 183434 75200
rect 249610 75148 249616 75200
rect 249668 75188 249674 75200
rect 546494 75188 546500 75200
rect 249668 75160 546500 75188
rect 249668 75148 249674 75160
rect 546494 75148 546500 75160
rect 546552 75148 546558 75200
rect 160002 75080 160008 75132
rect 160060 75120 160066 75132
rect 160278 75120 160284 75132
rect 160060 75092 160284 75120
rect 160060 75080 160066 75092
rect 160278 75080 160284 75092
rect 160336 75080 160342 75132
rect 179322 75080 179328 75132
rect 179380 75120 179386 75132
rect 179598 75120 179604 75132
rect 179380 75092 179604 75120
rect 179380 75080 179386 75092
rect 179598 75080 179604 75092
rect 179656 75080 179662 75132
rect 184842 75080 184848 75132
rect 184900 75120 184906 75132
rect 185118 75120 185124 75132
rect 184900 75092 185124 75120
rect 184900 75080 184906 75092
rect 185118 75080 185124 75092
rect 185176 75080 185182 75132
rect 160186 75012 160192 75064
rect 160244 75052 160250 75064
rect 160738 75052 160744 75064
rect 160244 75024 160744 75052
rect 160244 75012 160250 75024
rect 160738 75012 160744 75024
rect 160796 75012 160802 75064
rect 179506 75012 179512 75064
rect 179564 75052 179570 75064
rect 180058 75052 180064 75064
rect 179564 75024 180064 75052
rect 179564 75012 179570 75024
rect 180058 75012 180064 75024
rect 180116 75012 180122 75064
rect 185026 75012 185032 75064
rect 185084 75052 185090 75064
rect 185946 75052 185952 75064
rect 185084 75024 185952 75052
rect 185084 75012 185090 75024
rect 185946 75012 185952 75024
rect 186004 75012 186010 75064
rect 167454 74060 167460 74112
rect 167512 74100 167518 74112
rect 284294 74100 284300 74112
rect 167512 74072 284300 74100
rect 167512 74060 167518 74072
rect 284294 74060 284300 74072
rect 284352 74060 284358 74112
rect 212626 73992 212632 74044
rect 212684 74032 212690 74044
rect 431954 74032 431960 74044
rect 212684 74004 431960 74032
rect 212684 73992 212690 74004
rect 431954 73992 431960 74004
rect 432012 73992 432018 74044
rect 239030 73924 239036 73976
rect 239088 73964 239094 73976
rect 514754 73964 514760 73976
rect 239088 73936 514760 73964
rect 239088 73924 239094 73936
rect 514754 73924 514760 73936
rect 514812 73924 514818 73976
rect 243170 73856 243176 73908
rect 243228 73896 243234 73908
rect 527174 73896 527180 73908
rect 243228 73868 527180 73896
rect 243228 73856 243234 73868
rect 527174 73856 527180 73868
rect 527232 73856 527238 73908
rect 247310 73788 247316 73840
rect 247368 73828 247374 73840
rect 540974 73828 540980 73840
rect 247368 73800 540980 73828
rect 247368 73788 247374 73800
rect 540974 73788 540980 73800
rect 541032 73788 541038 73840
rect 561122 73108 561128 73160
rect 561180 73148 561186 73160
rect 579982 73148 579988 73160
rect 561180 73120 579988 73148
rect 561180 73108 561186 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 166626 72700 166632 72752
rect 166684 72740 166690 72752
rect 280154 72740 280160 72752
rect 166684 72712 280160 72740
rect 166684 72700 166690 72712
rect 280154 72700 280160 72712
rect 280212 72700 280218 72752
rect 196710 72632 196716 72684
rect 196768 72672 196774 72684
rect 378134 72672 378140 72684
rect 196768 72644 378140 72672
rect 196768 72632 196774 72644
rect 378134 72632 378140 72644
rect 378192 72632 378198 72684
rect 211798 72564 211804 72616
rect 211856 72604 211862 72616
rect 427814 72604 427820 72616
rect 211856 72576 427820 72604
rect 211856 72564 211862 72576
rect 427814 72564 427820 72576
rect 427872 72564 427878 72616
rect 243078 72496 243084 72548
rect 243136 72536 243142 72548
rect 529934 72536 529940 72548
rect 243136 72508 529940 72536
rect 243136 72496 243142 72508
rect 529934 72496 529940 72508
rect 529992 72496 529998 72548
rect 247218 72428 247224 72480
rect 247276 72468 247282 72480
rect 539594 72468 539600 72480
rect 247276 72440 539600 72468
rect 247276 72428 247282 72440
rect 539594 72428 539600 72440
rect 539652 72428 539658 72480
rect 165522 71272 165528 71324
rect 165580 71312 165586 71324
rect 276014 71312 276020 71324
rect 165580 71284 276020 71312
rect 165580 71272 165586 71284
rect 276014 71272 276020 71284
rect 276072 71272 276078 71324
rect 207106 71204 207112 71256
rect 207164 71244 207170 71256
rect 414014 71244 414020 71256
rect 207164 71216 414020 71244
rect 207164 71204 207170 71216
rect 414014 71204 414020 71216
rect 414072 71204 414078 71256
rect 209958 71136 209964 71188
rect 210016 71176 210022 71188
rect 420914 71176 420920 71188
rect 210016 71148 420920 71176
rect 210016 71136 210022 71148
rect 420914 71136 420920 71148
rect 420972 71136 420978 71188
rect 211338 71068 211344 71120
rect 211396 71108 211402 71120
rect 423674 71108 423680 71120
rect 211396 71080 423680 71108
rect 211396 71068 211402 71080
rect 423674 71068 423680 71080
rect 423732 71068 423738 71120
rect 255590 71000 255596 71052
rect 255648 71040 255654 71052
rect 571334 71040 571340 71052
rect 255648 71012 571340 71040
rect 255648 71000 255654 71012
rect 571334 71000 571340 71012
rect 571392 71000 571398 71052
rect 164418 69912 164424 69964
rect 164476 69952 164482 69964
rect 273254 69952 273260 69964
rect 164476 69924 273260 69952
rect 164476 69912 164482 69924
rect 273254 69912 273260 69924
rect 273312 69912 273318 69964
rect 197814 69844 197820 69896
rect 197872 69884 197878 69896
rect 382274 69884 382280 69896
rect 197872 69856 382280 69884
rect 197872 69844 197878 69856
rect 382274 69844 382280 69856
rect 382332 69844 382338 69896
rect 203426 69776 203432 69828
rect 203484 69816 203490 69828
rect 398834 69816 398840 69828
rect 203484 69788 398840 69816
rect 203484 69776 203490 69788
rect 398834 69776 398840 69788
rect 398892 69776 398898 69828
rect 204438 69708 204444 69760
rect 204496 69748 204502 69760
rect 402974 69748 402980 69760
rect 204496 69720 402980 69748
rect 204496 69708 204502 69720
rect 402974 69708 402980 69720
rect 403032 69708 403038 69760
rect 254210 69640 254216 69692
rect 254268 69680 254274 69692
rect 564526 69680 564532 69692
rect 254268 69652 564532 69680
rect 254268 69640 254274 69652
rect 564526 69640 564532 69652
rect 564584 69640 564590 69692
rect 163130 68552 163136 68604
rect 163188 68592 163194 68604
rect 269114 68592 269120 68604
rect 163188 68564 269120 68592
rect 163188 68552 163194 68564
rect 269114 68552 269120 68564
rect 269172 68552 269178 68604
rect 199010 68484 199016 68536
rect 199068 68524 199074 68536
rect 385034 68524 385040 68536
rect 199068 68496 385040 68524
rect 199068 68484 199074 68496
rect 385034 68484 385040 68496
rect 385092 68484 385098 68536
rect 200390 68416 200396 68468
rect 200448 68456 200454 68468
rect 391934 68456 391940 68468
rect 200448 68428 391940 68456
rect 200448 68416 200454 68428
rect 391934 68416 391940 68428
rect 391992 68416 391998 68468
rect 202138 68348 202144 68400
rect 202196 68388 202202 68400
rect 396074 68388 396080 68400
rect 202196 68360 396080 68388
rect 202196 68348 202202 68360
rect 396074 68348 396080 68360
rect 396132 68348 396138 68400
rect 251450 68280 251456 68332
rect 251508 68320 251514 68332
rect 556154 68320 556160 68332
rect 251508 68292 556160 68320
rect 251508 68280 251514 68292
rect 556154 68280 556160 68292
rect 556212 68280 556218 68332
rect 162026 67124 162032 67176
rect 162084 67164 162090 67176
rect 266354 67164 266360 67176
rect 162084 67136 266360 67164
rect 162084 67124 162090 67136
rect 266354 67124 266360 67136
rect 266412 67124 266418 67176
rect 189718 67056 189724 67108
rect 189776 67096 189782 67108
rect 357434 67096 357440 67108
rect 189776 67068 357440 67096
rect 189776 67056 189782 67068
rect 357434 67056 357440 67068
rect 357492 67056 357498 67108
rect 194778 66988 194784 67040
rect 194836 67028 194842 67040
rect 371234 67028 371240 67040
rect 194836 67000 371240 67028
rect 194836 66988 194842 67000
rect 371234 66988 371240 67000
rect 371292 66988 371298 67040
rect 200298 66920 200304 66972
rect 200356 66960 200362 66972
rect 389174 66960 389180 66972
rect 200356 66932 389180 66960
rect 200356 66920 200362 66932
rect 389174 66920 389180 66932
rect 389232 66920 389238 66972
rect 250438 66852 250444 66904
rect 250496 66892 250502 66904
rect 553394 66892 553400 66904
rect 250496 66864 553400 66892
rect 250496 66852 250502 66864
rect 553394 66852 553400 66864
rect 553452 66852 553458 66904
rect 160922 65764 160928 65816
rect 160980 65804 160986 65816
rect 262214 65804 262220 65816
rect 160980 65776 262220 65804
rect 160980 65764 160986 65776
rect 262214 65764 262220 65776
rect 262272 65764 262278 65816
rect 186866 65696 186872 65748
rect 186924 65736 186930 65748
rect 346394 65736 346400 65748
rect 186924 65708 346400 65736
rect 186924 65696 186930 65708
rect 346394 65696 346400 65708
rect 346452 65696 346458 65748
rect 187878 65628 187884 65680
rect 187936 65668 187942 65680
rect 349154 65668 349160 65680
rect 187936 65640 349160 65668
rect 187936 65628 187942 65640
rect 349154 65628 349160 65640
rect 349212 65628 349218 65680
rect 92750 65560 92756 65612
rect 92808 65560 92814 65612
rect 189166 65560 189172 65612
rect 189224 65600 189230 65612
rect 353294 65600 353300 65612
rect 189224 65572 353300 65600
rect 189224 65560 189230 65572
rect 353294 65560 353300 65572
rect 353352 65560 353358 65612
rect 92768 65408 92796 65560
rect 247126 65492 247132 65544
rect 247184 65532 247190 65544
rect 542354 65532 542360 65544
rect 247184 65504 542360 65532
rect 247184 65492 247190 65504
rect 542354 65492 542360 65504
rect 542412 65492 542418 65544
rect 92750 65356 92756 65408
rect 92808 65356 92814 65408
rect 160278 64404 160284 64456
rect 160336 64444 160342 64456
rect 259546 64444 259552 64456
rect 160336 64416 259552 64444
rect 160336 64404 160342 64416
rect 259546 64404 259552 64416
rect 259604 64404 259610 64456
rect 183738 64336 183744 64388
rect 183796 64376 183802 64388
rect 335354 64376 335360 64388
rect 183796 64348 335360 64376
rect 183796 64336 183802 64348
rect 335354 64336 335360 64348
rect 335412 64336 335418 64388
rect 185118 64268 185124 64320
rect 185176 64308 185182 64320
rect 339494 64308 339500 64320
rect 185176 64280 339500 64308
rect 185176 64268 185182 64280
rect 339494 64268 339500 64280
rect 339552 64268 339558 64320
rect 185026 64200 185032 64252
rect 185084 64240 185090 64252
rect 342254 64240 342260 64252
rect 185084 64212 342260 64240
rect 185084 64200 185090 64212
rect 342254 64200 342260 64212
rect 342312 64200 342318 64252
rect 238938 64132 238944 64184
rect 238996 64172 239002 64184
rect 517514 64172 517520 64184
rect 238996 64144 517520 64172
rect 238996 64132 239002 64144
rect 517514 64132 517520 64144
rect 517572 64132 517578 64184
rect 169938 63044 169944 63096
rect 169996 63084 170002 63096
rect 293954 63084 293960 63096
rect 169996 63056 293960 63084
rect 169996 63044 170002 63056
rect 293954 63044 293960 63056
rect 294012 63044 294018 63096
rect 179690 62976 179696 63028
rect 179748 63016 179754 63028
rect 324314 63016 324320 63028
rect 179748 62988 324320 63016
rect 179748 62976 179754 62988
rect 324314 62976 324320 62988
rect 324372 62976 324378 63028
rect 181070 62908 181076 62960
rect 181128 62948 181134 62960
rect 328454 62948 328460 62960
rect 181128 62920 328460 62948
rect 181128 62908 181134 62920
rect 328454 62908 328460 62920
rect 328512 62908 328518 62960
rect 182450 62840 182456 62892
rect 182508 62880 182514 62892
rect 332594 62880 332600 62892
rect 182508 62852 332600 62880
rect 182508 62840 182514 62852
rect 332594 62840 332600 62852
rect 332652 62840 332658 62892
rect 117314 62772 117320 62824
rect 117372 62812 117378 62824
rect 117498 62812 117504 62824
rect 117372 62784 117504 62812
rect 117372 62772 117378 62784
rect 117498 62772 117504 62784
rect 117556 62772 117562 62824
rect 238846 62772 238852 62824
rect 238904 62812 238910 62824
rect 514846 62812 514852 62824
rect 238904 62784 514852 62812
rect 238904 62772 238910 62784
rect 514846 62772 514852 62784
rect 514904 62772 514910 62824
rect 176930 61616 176936 61668
rect 176988 61656 176994 61668
rect 314654 61656 314660 61668
rect 176988 61628 314660 61656
rect 176988 61616 176994 61628
rect 314654 61616 314660 61628
rect 314712 61616 314718 61668
rect 178126 61548 178132 61600
rect 178184 61588 178190 61600
rect 317414 61588 317420 61600
rect 178184 61560 317420 61588
rect 178184 61548 178190 61560
rect 317414 61548 317420 61560
rect 317472 61548 317478 61600
rect 179598 61480 179604 61532
rect 179656 61520 179662 61532
rect 321554 61520 321560 61532
rect 179656 61492 321560 61520
rect 179656 61480 179662 61492
rect 321554 61480 321560 61492
rect 321612 61480 321618 61532
rect 194686 61412 194692 61464
rect 194744 61452 194750 61464
rect 372614 61452 372620 61464
rect 194744 61424 372620 61452
rect 194744 61412 194750 61424
rect 372614 61412 372620 61424
rect 372672 61412 372678 61464
rect 229370 61344 229376 61396
rect 229428 61384 229434 61396
rect 485774 61384 485780 61396
rect 229428 61356 485780 61384
rect 229428 61344 229434 61356
rect 485774 61344 485780 61356
rect 485832 61344 485838 61396
rect 561030 60664 561036 60716
rect 561088 60704 561094 60716
rect 580166 60704 580172 60716
rect 561088 60676 580172 60704
rect 561088 60664 561094 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 174078 60256 174084 60308
rect 174136 60296 174142 60308
rect 303614 60296 303620 60308
rect 174136 60268 303620 60296
rect 174136 60256 174142 60268
rect 303614 60256 303620 60268
rect 303672 60256 303678 60308
rect 174170 60188 174176 60240
rect 174228 60228 174234 60240
rect 307754 60228 307760 60240
rect 174228 60200 307760 60228
rect 174228 60188 174234 60200
rect 307754 60188 307760 60200
rect 307812 60188 307818 60240
rect 175550 60120 175556 60172
rect 175608 60160 175614 60172
rect 310514 60160 310520 60172
rect 175608 60132 310520 60160
rect 175608 60120 175614 60132
rect 310514 60120 310520 60132
rect 310572 60120 310578 60172
rect 247034 60052 247040 60104
rect 247092 60092 247098 60104
rect 543734 60092 543740 60104
rect 247092 60064 543740 60092
rect 247092 60052 247098 60064
rect 543734 60052 543740 60064
rect 543792 60052 543798 60104
rect 149146 59984 149152 60036
rect 149204 60024 149210 60036
rect 223666 60024 223672 60036
rect 149204 59996 223672 60024
rect 149204 59984 149210 59996
rect 223666 59984 223672 59996
rect 223724 59984 223730 60036
rect 258166 59984 258172 60036
rect 258224 60024 258230 60036
rect 576854 60024 576860 60036
rect 258224 59996 576860 60024
rect 258224 59984 258230 59996
rect 576854 59984 576860 59996
rect 576912 59984 576918 60036
rect 169846 58964 169852 59016
rect 169904 59004 169910 59016
rect 292574 59004 292580 59016
rect 169904 58976 292580 59004
rect 169904 58964 169910 58976
rect 292574 58964 292580 58976
rect 292632 58964 292638 59016
rect 171318 58896 171324 58948
rect 171376 58936 171382 58948
rect 296714 58936 296720 58948
rect 171376 58908 296720 58936
rect 171376 58896 171382 58908
rect 296714 58896 296720 58908
rect 296772 58896 296778 58948
rect 225138 58828 225144 58880
rect 225196 58868 225202 58880
rect 471974 58868 471980 58880
rect 225196 58840 471980 58868
rect 225196 58828 225202 58840
rect 471974 58828 471980 58840
rect 472032 58828 472038 58880
rect 253934 58760 253940 58812
rect 253992 58800 253998 58812
rect 563054 58800 563060 58812
rect 253992 58772 563060 58800
rect 253992 58760 253998 58772
rect 563054 58760 563060 58772
rect 563112 58760 563118 58812
rect 254118 58692 254124 58744
rect 254176 58732 254182 58744
rect 565814 58732 565820 58744
rect 254176 58704 565820 58732
rect 254176 58692 254182 58704
rect 565814 58692 565820 58704
rect 565872 58692 565878 58744
rect 255498 58624 255504 58676
rect 255556 58664 255562 58676
rect 569954 58664 569960 58676
rect 255556 58636 569960 58664
rect 255556 58624 255562 58636
rect 569954 58624 569960 58636
rect 570012 58624 570018 58676
rect 92658 58556 92664 58608
rect 92716 58596 92722 58608
rect 92842 58596 92848 58608
rect 92716 58568 92848 58596
rect 92716 58556 92722 58568
rect 92842 58556 92848 58568
rect 92900 58556 92906 58608
rect 168558 57536 168564 57588
rect 168616 57576 168622 57588
rect 285674 57576 285680 57588
rect 168616 57548 285680 57576
rect 168616 57536 168622 57548
rect 285674 57536 285680 57548
rect 285732 57536 285738 57588
rect 168466 57468 168472 57520
rect 168524 57508 168530 57520
rect 289814 57508 289820 57520
rect 168524 57480 289820 57508
rect 168524 57468 168530 57480
rect 289814 57468 289820 57480
rect 289872 57468 289878 57520
rect 223850 57400 223856 57452
rect 223908 57440 223914 57452
rect 465074 57440 465080 57452
rect 223908 57412 465080 57440
rect 223908 57400 223914 57412
rect 465074 57400 465080 57412
rect 465132 57400 465138 57452
rect 244550 57332 244556 57384
rect 244608 57372 244614 57384
rect 534074 57372 534080 57384
rect 244608 57344 534080 57372
rect 244608 57332 244614 57344
rect 534074 57332 534080 57344
rect 534132 57332 534138 57384
rect 245838 57264 245844 57316
rect 245896 57304 245902 57316
rect 538214 57304 538220 57316
rect 245896 57276 538220 57304
rect 245896 57264 245902 57276
rect 538214 57264 538220 57276
rect 538272 57264 538278 57316
rect 248598 57196 248604 57248
rect 248656 57236 248662 57248
rect 545114 57236 545120 57248
rect 248656 57208 545120 57236
rect 248656 57196 248662 57208
rect 545114 57196 545120 57208
rect 545172 57196 545178 57248
rect 165706 56176 165712 56228
rect 165764 56216 165770 56228
rect 278774 56216 278780 56228
rect 165764 56188 278780 56216
rect 165764 56176 165770 56188
rect 278774 56176 278780 56188
rect 278832 56176 278838 56228
rect 167086 56108 167092 56160
rect 167144 56148 167150 56160
rect 282914 56148 282920 56160
rect 167144 56120 282920 56148
rect 167144 56108 167150 56120
rect 282914 56108 282920 56120
rect 282972 56108 282978 56160
rect 220998 56040 221004 56092
rect 221056 56080 221062 56092
rect 456794 56080 456800 56092
rect 221056 56052 456800 56080
rect 221056 56040 221062 56052
rect 456794 56040 456800 56052
rect 456852 56040 456858 56092
rect 240318 55972 240324 56024
rect 240376 56012 240382 56024
rect 520274 56012 520280 56024
rect 240376 55984 520280 56012
rect 240376 55972 240382 55984
rect 520274 55972 520280 55984
rect 520332 55972 520338 56024
rect 241790 55904 241796 55956
rect 241848 55944 241854 55956
rect 523034 55944 523040 55956
rect 241848 55916 523040 55944
rect 241848 55904 241854 55916
rect 523034 55904 523040 55916
rect 523092 55904 523098 55956
rect 242986 55836 242992 55888
rect 243044 55876 243050 55888
rect 531314 55876 531320 55888
rect 243044 55848 531320 55876
rect 243044 55836 243050 55848
rect 531314 55836 531320 55848
rect 531372 55836 531378 55888
rect 164326 54816 164332 54868
rect 164384 54856 164390 54868
rect 276106 54856 276112 54868
rect 164384 54828 276112 54856
rect 164384 54816 164390 54828
rect 276106 54816 276112 54828
rect 276164 54816 276170 54868
rect 218330 54748 218336 54800
rect 218388 54788 218394 54800
rect 447134 54788 447140 54800
rect 218388 54760 447140 54788
rect 218388 54748 218394 54760
rect 447134 54748 447140 54760
rect 447192 54748 447198 54800
rect 237466 54680 237472 54732
rect 237524 54720 237530 54732
rect 509234 54720 509240 54732
rect 237524 54692 509240 54720
rect 237524 54680 237530 54692
rect 509234 54680 509240 54692
rect 509292 54680 509298 54732
rect 237650 54612 237656 54664
rect 237708 54652 237714 54664
rect 513374 54652 513380 54664
rect 237708 54624 513380 54652
rect 237708 54612 237714 54624
rect 513374 54612 513380 54624
rect 513432 54612 513438 54664
rect 238754 54544 238760 54596
rect 238812 54584 238818 54596
rect 516134 54584 516140 54596
rect 238812 54556 516140 54584
rect 238812 54544 238818 54556
rect 516134 54544 516140 54556
rect 516192 54544 516198 54596
rect 256878 54476 256884 54528
rect 256936 54516 256942 54528
rect 572714 54516 572720 54528
rect 256936 54488 572720 54516
rect 256936 54476 256942 54488
rect 572714 54476 572720 54488
rect 572772 54476 572778 54528
rect 163038 53388 163044 53440
rect 163096 53428 163102 53440
rect 267734 53428 267740 53440
rect 163096 53400 267740 53428
rect 163096 53388 163102 53400
rect 267734 53388 267740 53400
rect 267792 53388 267798 53440
rect 162946 53320 162952 53372
rect 163004 53360 163010 53372
rect 271874 53360 271880 53372
rect 163004 53332 271880 53360
rect 163004 53320 163010 53332
rect 271874 53320 271880 53332
rect 271932 53320 271938 53372
rect 214098 53252 214104 53304
rect 214156 53292 214162 53304
rect 436094 53292 436100 53304
rect 214156 53264 436100 53292
rect 214156 53252 214162 53264
rect 436094 53252 436100 53264
rect 436152 53252 436158 53304
rect 233418 53184 233424 53236
rect 233476 53224 233482 53236
rect 498194 53224 498200 53236
rect 233476 53196 498200 53224
rect 233476 53184 233482 53196
rect 498194 53184 498200 53196
rect 498252 53184 498258 53236
rect 234890 53116 234896 53168
rect 234948 53156 234954 53168
rect 502334 53156 502340 53168
rect 234948 53128 502340 53156
rect 234948 53116 234954 53128
rect 502334 53116 502340 53128
rect 502392 53116 502398 53168
rect 236270 53048 236276 53100
rect 236328 53088 236334 53100
rect 506474 53088 506480 53100
rect 236328 53060 506480 53088
rect 236328 53048 236334 53060
rect 506474 53048 506480 53060
rect 506532 53048 506538 53100
rect 153286 52028 153292 52080
rect 153344 52068 153350 52080
rect 237466 52068 237472 52080
rect 153344 52040 237472 52068
rect 153344 52028 153350 52040
rect 237466 52028 237472 52040
rect 237524 52028 237530 52080
rect 161658 51960 161664 52012
rect 161716 52000 161722 52012
rect 264974 52000 264980 52012
rect 161716 51972 264980 52000
rect 161716 51960 161722 51972
rect 264974 51960 264980 51972
rect 265032 51960 265038 52012
rect 171226 51892 171232 51944
rect 171284 51932 171290 51944
rect 298094 51932 298100 51944
rect 171284 51904 298100 51932
rect 171284 51892 171290 51904
rect 298094 51892 298100 51904
rect 298152 51892 298158 51944
rect 226518 51824 226524 51876
rect 226576 51864 226582 51876
rect 476114 51864 476120 51876
rect 226576 51836 476120 51864
rect 226576 51824 226582 51836
rect 476114 51824 476120 51836
rect 476172 51824 476178 51876
rect 232038 51756 232044 51808
rect 232096 51796 232102 51808
rect 491294 51796 491300 51808
rect 232096 51768 491300 51796
rect 232096 51756 232102 51768
rect 491294 51756 491300 51768
rect 491352 51756 491358 51808
rect 232130 51688 232136 51740
rect 232188 51728 232194 51740
rect 495434 51728 495440 51740
rect 232188 51700 495440 51728
rect 232188 51688 232194 51700
rect 495434 51688 495440 51700
rect 495492 51688 495498 51740
rect 152090 50668 152096 50720
rect 152148 50708 152154 50720
rect 234890 50708 234896 50720
rect 152148 50680 234896 50708
rect 152148 50668 152154 50680
rect 234890 50668 234896 50680
rect 234948 50668 234954 50720
rect 160186 50600 160192 50652
rect 160244 50640 160250 50652
rect 260834 50640 260840 50652
rect 160244 50612 260840 50640
rect 160244 50600 160250 50612
rect 260834 50600 260840 50612
rect 260892 50600 260898 50652
rect 195238 50532 195244 50584
rect 195296 50572 195302 50584
rect 368474 50572 368480 50584
rect 195296 50544 368480 50572
rect 195296 50532 195302 50544
rect 368474 50532 368480 50544
rect 368532 50532 368538 50584
rect 222378 50464 222384 50516
rect 222436 50504 222442 50516
rect 462314 50504 462320 50516
rect 222436 50476 462320 50504
rect 222436 50464 222442 50476
rect 462314 50464 462320 50476
rect 462372 50464 462378 50516
rect 223758 50396 223764 50448
rect 223816 50436 223822 50448
rect 465166 50436 465172 50448
rect 223816 50408 465172 50436
rect 223816 50396 223822 50408
rect 465166 50396 465172 50408
rect 465224 50396 465230 50448
rect 137278 50328 137284 50380
rect 137336 50368 137342 50380
rect 178126 50368 178132 50380
rect 137336 50340 178132 50368
rect 137336 50328 137342 50340
rect 178126 50328 178132 50340
rect 178184 50328 178190 50380
rect 225046 50328 225052 50380
rect 225104 50368 225110 50380
rect 473354 50368 473360 50380
rect 225104 50340 473360 50368
rect 225104 50328 225110 50340
rect 473354 50328 473360 50340
rect 473412 50328 473418 50380
rect 158898 49240 158904 49292
rect 158956 49280 158962 49292
rect 258166 49280 258172 49292
rect 158956 49252 258172 49280
rect 158956 49240 158962 49252
rect 258166 49240 258172 49252
rect 258224 49240 258230 49292
rect 191282 49172 191288 49224
rect 191340 49212 191346 49224
rect 354674 49212 354680 49224
rect 191340 49184 354680 49212
rect 191340 49172 191346 49184
rect 354674 49172 354680 49184
rect 354732 49172 354738 49224
rect 219618 49104 219624 49156
rect 219676 49144 219682 49156
rect 451274 49144 451280 49156
rect 219676 49116 451280 49144
rect 219676 49104 219682 49116
rect 451274 49104 451280 49116
rect 451332 49104 451338 49156
rect 219526 49036 219532 49088
rect 219584 49076 219590 49088
rect 455414 49076 455420 49088
rect 219584 49048 455420 49076
rect 219584 49036 219590 49048
rect 455414 49036 455420 49048
rect 455472 49036 455478 49088
rect 52454 48968 52460 49020
rect 52512 49008 52518 49020
rect 95418 49008 95424 49020
rect 52512 48980 95424 49008
rect 52512 48968 52518 48980
rect 95418 48968 95424 48980
rect 95476 48968 95482 49020
rect 220906 48968 220912 49020
rect 220964 49008 220970 49020
rect 458174 49008 458180 49020
rect 220964 48980 458180 49008
rect 220964 48968 220970 48980
rect 458174 48968 458180 48980
rect 458232 48968 458238 49020
rect 157610 47880 157616 47932
rect 157668 47920 157674 47932
rect 253934 47920 253940 47932
rect 157668 47892 253940 47920
rect 157668 47880 157674 47892
rect 253934 47880 253940 47892
rect 253992 47880 253998 47932
rect 226978 47812 226984 47864
rect 227036 47852 227042 47864
rect 440326 47852 440332 47864
rect 227036 47824 440332 47852
rect 227036 47812 227042 47824
rect 440326 47812 440332 47824
rect 440384 47812 440390 47864
rect 215294 47744 215300 47796
rect 215352 47784 215358 47796
rect 440234 47784 440240 47796
rect 215352 47756 440240 47784
rect 215352 47744 215358 47756
rect 440234 47744 440240 47756
rect 440292 47744 440298 47796
rect 216766 47676 216772 47728
rect 216824 47716 216830 47728
rect 444374 47716 444380 47728
rect 216824 47688 444380 47716
rect 216824 47676 216830 47688
rect 444374 47676 444380 47688
rect 444432 47676 444438 47728
rect 218238 47608 218244 47660
rect 218296 47648 218302 47660
rect 448514 47648 448520 47660
rect 218296 47620 448520 47648
rect 218296 47608 218302 47620
rect 448514 47608 448520 47620
rect 448572 47608 448578 47660
rect 147950 47540 147956 47592
rect 148008 47580 148014 47592
rect 219526 47580 219532 47592
rect 148008 47552 219532 47580
rect 148008 47540 148014 47552
rect 219526 47540 219532 47552
rect 219584 47540 219590 47592
rect 244458 47540 244464 47592
rect 244516 47580 244522 47592
rect 535454 47580 535460 47592
rect 244516 47552 535460 47580
rect 244516 47540 244522 47552
rect 535454 47540 535460 47552
rect 535512 47540 535518 47592
rect 261478 46860 261484 46912
rect 261536 46900 261542 46912
rect 550082 46900 550088 46912
rect 261536 46872 550088 46900
rect 261536 46860 261542 46872
rect 550082 46860 550088 46872
rect 550140 46900 550146 46912
rect 550542 46900 550548 46912
rect 550140 46872 550548 46900
rect 550140 46860 550146 46872
rect 550542 46860 550548 46872
rect 550600 46860 550606 46912
rect 157518 46452 157524 46504
rect 157576 46492 157582 46504
rect 251450 46492 251456 46504
rect 157576 46464 251456 46492
rect 157576 46452 157582 46464
rect 251450 46452 251456 46464
rect 251508 46452 251514 46504
rect 192018 46384 192024 46436
rect 192076 46424 192082 46436
rect 361574 46424 361580 46436
rect 192076 46396 361580 46424
rect 192076 46384 192082 46396
rect 361574 46384 361580 46396
rect 361632 46384 361638 46436
rect 196066 46316 196072 46368
rect 196124 46356 196130 46368
rect 376754 46356 376760 46368
rect 196124 46328 376760 46356
rect 196124 46316 196130 46328
rect 376754 46316 376760 46328
rect 376812 46316 376818 46368
rect 204346 46248 204352 46300
rect 204404 46288 204410 46300
rect 405734 46288 405740 46300
rect 204404 46260 405740 46288
rect 204404 46248 204410 46260
rect 405734 46248 405740 46260
rect 405792 46248 405798 46300
rect 207014 46180 207020 46232
rect 207072 46220 207078 46232
rect 412634 46220 412640 46232
rect 207072 46192 412640 46220
rect 207072 46180 207078 46192
rect 412634 46180 412640 46192
rect 412692 46180 412698 46232
rect 550542 46180 550548 46232
rect 550600 46220 550606 46232
rect 580166 46220 580172 46232
rect 550600 46192 580172 46220
rect 550600 46180 550606 46192
rect 580166 46180 580172 46192
rect 580224 46180 580230 46232
rect 169018 45092 169024 45144
rect 169076 45132 169082 45144
rect 281534 45132 281540 45144
rect 169076 45104 281540 45132
rect 169076 45092 169082 45104
rect 281534 45092 281540 45104
rect 281592 45092 281598 45144
rect 189074 45024 189080 45076
rect 189132 45064 189138 45076
rect 356054 45064 356060 45076
rect 189132 45036 356060 45064
rect 189132 45024 189138 45036
rect 356054 45024 356060 45036
rect 356112 45024 356118 45076
rect 193398 44956 193404 45008
rect 193456 44996 193462 45008
rect 369854 44996 369860 45008
rect 193456 44968 369860 44996
rect 193456 44956 193462 44968
rect 369854 44956 369860 44968
rect 369912 44956 369918 45008
rect 138290 44888 138296 44940
rect 138348 44928 138354 44940
rect 184198 44928 184204 44940
rect 138348 44900 184204 44928
rect 138348 44888 138354 44900
rect 184198 44888 184204 44900
rect 184256 44888 184262 44940
rect 211246 44888 211252 44940
rect 211304 44928 211310 44940
rect 425054 44928 425060 44940
rect 211304 44900 425060 44928
rect 211304 44888 211310 44900
rect 425054 44888 425060 44900
rect 425112 44888 425118 44940
rect 30374 44820 30380 44872
rect 30432 44860 30438 44872
rect 88518 44860 88524 44872
rect 30432 44832 88524 44860
rect 30432 44820 30438 44832
rect 88518 44820 88524 44832
rect 88576 44820 88582 44872
rect 145190 44820 145196 44872
rect 145248 44860 145254 44872
rect 210510 44860 210516 44872
rect 145248 44832 210516 44860
rect 145248 44820 145254 44832
rect 210510 44820 210516 44832
rect 210568 44820 210574 44872
rect 229278 44820 229284 44872
rect 229336 44860 229342 44872
rect 481634 44860 481640 44872
rect 229336 44832 481640 44860
rect 229336 44820 229342 44832
rect 481634 44820 481640 44832
rect 481692 44820 481698 44872
rect 156230 43732 156236 43784
rect 156288 43772 156294 43784
rect 247034 43772 247040 43784
rect 156288 43744 247040 43772
rect 156288 43732 156294 43744
rect 247034 43732 247040 43744
rect 247092 43732 247098 43784
rect 211154 43664 211160 43716
rect 211212 43704 211218 43716
rect 426434 43704 426440 43716
rect 211212 43676 426440 43704
rect 211212 43664 211218 43676
rect 426434 43664 426440 43676
rect 426492 43664 426498 43716
rect 73154 43596 73160 43648
rect 73212 43636 73218 43648
rect 102318 43636 102324 43648
rect 73212 43608 102324 43636
rect 73212 43596 73218 43608
rect 102318 43596 102324 43608
rect 102376 43596 102382 43648
rect 215938 43596 215944 43648
rect 215996 43636 216002 43648
rect 432046 43636 432052 43648
rect 215996 43608 432052 43636
rect 215996 43596 216002 43608
rect 432046 43596 432052 43608
rect 432104 43596 432110 43648
rect 66254 43528 66260 43580
rect 66312 43568 66318 43580
rect 99558 43568 99564 43580
rect 66312 43540 99564 43568
rect 66312 43528 66318 43540
rect 99558 43528 99564 43540
rect 99616 43528 99622 43580
rect 212718 43528 212724 43580
rect 212776 43568 212782 43580
rect 430574 43568 430580 43580
rect 212776 43540 430580 43568
rect 212776 43528 212782 43540
rect 430574 43528 430580 43540
rect 430632 43528 430638 43580
rect 59354 43460 59360 43512
rect 59412 43500 59418 43512
rect 98270 43500 98276 43512
rect 59412 43472 98276 43500
rect 59412 43460 59418 43472
rect 98270 43460 98276 43472
rect 98328 43460 98334 43512
rect 214006 43460 214012 43512
rect 214064 43500 214070 43512
rect 433334 43500 433340 43512
rect 214064 43472 433340 43500
rect 214064 43460 214070 43472
rect 433334 43460 433340 43472
rect 433392 43460 433398 43512
rect 22094 43392 22100 43444
rect 22152 43432 22158 43444
rect 87230 43432 87236 43444
rect 22152 43404 87236 43432
rect 22152 43392 22158 43404
rect 87230 43392 87236 43404
rect 87288 43392 87294 43444
rect 102318 43392 102324 43444
rect 102376 43432 102382 43444
rect 110690 43432 110696 43444
rect 102376 43404 110696 43432
rect 102376 43392 102382 43404
rect 110690 43392 110696 43404
rect 110748 43392 110754 43444
rect 145098 43392 145104 43444
rect 145156 43432 145162 43444
rect 212626 43432 212632 43444
rect 145156 43404 212632 43432
rect 145156 43392 145162 43404
rect 212626 43392 212632 43404
rect 212684 43392 212690 43444
rect 236178 43392 236184 43444
rect 236236 43432 236242 43444
rect 505094 43432 505100 43444
rect 236236 43404 505100 43432
rect 236236 43392 236242 43404
rect 505094 43392 505100 43404
rect 505152 43392 505158 43444
rect 171134 42304 171140 42356
rect 171192 42344 171198 42356
rect 295334 42344 295340 42356
rect 171192 42316 295340 42344
rect 171192 42304 171198 42316
rect 295334 42304 295340 42316
rect 295392 42304 295398 42356
rect 193858 42236 193864 42288
rect 193916 42276 193922 42288
rect 365714 42276 365720 42288
rect 193916 42248 365720 42276
rect 193916 42236 193922 42248
rect 365714 42236 365720 42248
rect 365772 42236 365778 42288
rect 35894 42168 35900 42220
rect 35952 42208 35958 42220
rect 91186 42208 91192 42220
rect 35952 42180 91192 42208
rect 35952 42168 35958 42180
rect 91186 42168 91192 42180
rect 91244 42168 91250 42220
rect 208486 42168 208492 42220
rect 208544 42208 208550 42220
rect 415394 42208 415400 42220
rect 208544 42180 415400 42208
rect 208544 42168 208550 42180
rect 415394 42168 415400 42180
rect 415452 42168 415458 42220
rect 16574 42100 16580 42152
rect 16632 42140 16638 42152
rect 84378 42140 84384 42152
rect 16632 42112 84384 42140
rect 16632 42100 16638 42112
rect 84378 42100 84384 42112
rect 84436 42100 84442 42152
rect 209866 42100 209872 42152
rect 209924 42140 209930 42152
rect 419534 42140 419540 42152
rect 209924 42112 419540 42140
rect 209924 42100 209930 42112
rect 419534 42100 419540 42112
rect 419592 42100 419598 42152
rect 1394 42032 1400 42084
rect 1452 42072 1458 42084
rect 80330 42072 80336 42084
rect 1452 42044 80336 42072
rect 1452 42032 1458 42044
rect 80330 42032 80336 42044
rect 80388 42032 80394 42084
rect 125870 42032 125876 42084
rect 125928 42072 125934 42084
rect 149146 42072 149152 42084
rect 125928 42044 149152 42072
rect 125928 42032 125934 42044
rect 149146 42032 149152 42044
rect 149204 42032 149210 42084
rect 149238 42032 149244 42084
rect 149296 42072 149302 42084
rect 226518 42072 226524 42084
rect 149296 42044 226524 42072
rect 149296 42032 149302 42044
rect 226518 42032 226524 42044
rect 226576 42032 226582 42084
rect 229186 42032 229192 42084
rect 229244 42072 229250 42084
rect 483014 42072 483020 42084
rect 229244 42044 483020 42072
rect 229244 42032 229250 42044
rect 483014 42032 483020 42044
rect 483072 42032 483078 42084
rect 162854 41012 162860 41064
rect 162912 41052 162918 41064
rect 270494 41052 270500 41064
rect 162912 41024 270500 41052
rect 162912 41012 162918 41024
rect 270494 41012 270500 41024
rect 270552 41012 270558 41064
rect 166994 40944 167000 40996
rect 167052 40984 167058 40996
rect 284386 40984 284392 40996
rect 167052 40956 284392 40984
rect 167052 40944 167058 40956
rect 284386 40944 284392 40956
rect 284444 40944 284450 40996
rect 94222 40876 94228 40928
rect 94280 40916 94286 40928
rect 109126 40916 109132 40928
rect 94280 40888 109132 40916
rect 94280 40876 94286 40888
rect 109126 40876 109132 40888
rect 109184 40876 109190 40928
rect 202874 40876 202880 40928
rect 202932 40916 202938 40928
rect 398926 40916 398932 40928
rect 202932 40888 398932 40916
rect 202932 40876 202938 40888
rect 398926 40876 398932 40888
rect 398984 40876 398990 40928
rect 129182 40808 129188 40860
rect 129240 40848 129246 40860
rect 154850 40848 154856 40860
rect 129240 40820 154856 40848
rect 129240 40808 129246 40820
rect 154850 40808 154856 40820
rect 154908 40808 154914 40860
rect 216674 40808 216680 40860
rect 216732 40848 216738 40860
rect 442994 40848 443000 40860
rect 216732 40820 443000 40848
rect 216732 40808 216738 40820
rect 442994 40808 443000 40820
rect 443052 40808 443058 40860
rect 44174 40740 44180 40792
rect 44232 40780 44238 40792
rect 94130 40780 94136 40792
rect 44232 40752 94136 40780
rect 44232 40740 44238 40752
rect 94130 40740 94136 40752
rect 94188 40740 94194 40792
rect 135254 40740 135260 40792
rect 135312 40780 135318 40792
rect 181070 40780 181076 40792
rect 135312 40752 181076 40780
rect 135312 40740 135318 40752
rect 181070 40740 181076 40752
rect 181128 40740 181134 40792
rect 242894 40740 242900 40792
rect 242952 40780 242958 40792
rect 528554 40780 528560 40792
rect 242952 40752 528560 40780
rect 242952 40740 242958 40752
rect 528554 40740 528560 40752
rect 528612 40740 528618 40792
rect 14 40672 20 40724
rect 72 40712 78 40724
rect 80238 40712 80244 40724
rect 72 40684 80244 40712
rect 72 40672 78 40684
rect 80238 40672 80244 40684
rect 80296 40672 80302 40724
rect 145006 40672 145012 40724
rect 145064 40712 145070 40724
rect 209866 40712 209872 40724
rect 145064 40684 209872 40712
rect 145064 40672 145070 40684
rect 209866 40672 209872 40684
rect 209924 40672 209930 40724
rect 252738 40672 252744 40724
rect 252796 40712 252802 40724
rect 559006 40712 559012 40724
rect 252796 40684 559012 40712
rect 252796 40672 252802 40684
rect 559006 40672 559012 40684
rect 559064 40672 559070 40724
rect 198918 39584 198924 39636
rect 198976 39624 198982 39636
rect 387794 39624 387800 39636
rect 198976 39596 387800 39624
rect 198976 39584 198982 39596
rect 387794 39584 387800 39596
rect 387852 39584 387858 39636
rect 200206 39516 200212 39568
rect 200264 39556 200270 39568
rect 390554 39556 390560 39568
rect 200264 39528 390560 39556
rect 200264 39516 200270 39528
rect 390554 39516 390560 39528
rect 390612 39516 390618 39568
rect 206278 39448 206284 39500
rect 206336 39488 206342 39500
rect 400214 39488 400220 39500
rect 206336 39460 400220 39488
rect 206336 39448 206342 39460
rect 400214 39448 400220 39460
rect 400272 39448 400278 39500
rect 204254 39380 204260 39432
rect 204312 39420 204318 39432
rect 401594 39420 401600 39432
rect 204312 39392 401600 39420
rect 204312 39380 204318 39392
rect 401594 39380 401600 39392
rect 401652 39380 401658 39432
rect 154942 39312 154948 39364
rect 155000 39352 155006 39364
rect 242894 39352 242900 39364
rect 155000 39324 242900 39352
rect 155000 39312 155006 39324
rect 242894 39312 242900 39324
rect 242952 39312 242958 39364
rect 244366 39312 244372 39364
rect 244424 39352 244430 39364
rect 531406 39352 531412 39364
rect 244424 39324 531412 39352
rect 244424 39312 244430 39324
rect 531406 39312 531412 39324
rect 531464 39312 531470 39364
rect 153194 38224 153200 38276
rect 153252 38264 153258 38276
rect 240318 38264 240324 38276
rect 153252 38236 240324 38264
rect 153252 38224 153258 38236
rect 240318 38224 240324 38236
rect 240376 38224 240382 38276
rect 194594 38156 194600 38208
rect 194652 38196 194658 38208
rect 374086 38196 374092 38208
rect 194652 38168 374092 38196
rect 194652 38156 194658 38168
rect 374086 38156 374092 38168
rect 374144 38156 374150 38208
rect 197446 38088 197452 38140
rect 197504 38128 197510 38140
rect 380894 38128 380900 38140
rect 197504 38100 380900 38128
rect 197504 38088 197510 38100
rect 380894 38088 380900 38100
rect 380952 38088 380958 38140
rect 198826 38020 198832 38072
rect 198884 38060 198890 38072
rect 383654 38060 383660 38072
rect 198884 38032 383660 38060
rect 198884 38020 198890 38032
rect 383654 38020 383660 38032
rect 383712 38020 383718 38072
rect 217318 37952 217324 38004
rect 217376 37992 217382 38004
rect 422294 37992 422300 38004
rect 217376 37964 422300 37992
rect 217376 37952 217382 37964
rect 422294 37952 422300 37964
rect 422352 37952 422358 38004
rect 237558 37884 237564 37936
rect 237616 37924 237622 37936
rect 510614 37924 510620 37936
rect 237616 37896 510620 37924
rect 237616 37884 237622 37896
rect 510614 37884 510620 37896
rect 510672 37884 510678 37936
rect 151998 36864 152004 36916
rect 152056 36904 152062 36916
rect 236178 36904 236184 36916
rect 152056 36876 236184 36904
rect 152056 36864 152062 36876
rect 236178 36864 236184 36876
rect 236236 36864 236242 36916
rect 186406 36796 186412 36848
rect 186464 36836 186470 36848
rect 345014 36836 345020 36848
rect 186464 36808 345020 36836
rect 186464 36796 186470 36808
rect 345014 36796 345020 36808
rect 345072 36796 345078 36848
rect 191926 36728 191932 36780
rect 191984 36768 191990 36780
rect 362954 36768 362960 36780
rect 191984 36740 362960 36768
rect 191984 36728 191990 36740
rect 362954 36728 362960 36740
rect 363012 36728 363018 36780
rect 193306 36660 193312 36712
rect 193364 36700 193370 36712
rect 365806 36700 365812 36712
rect 193364 36672 365812 36700
rect 193364 36660 193370 36672
rect 365806 36660 365812 36672
rect 365864 36660 365870 36712
rect 214558 36592 214564 36644
rect 214616 36632 214622 36644
rect 418154 36632 418160 36644
rect 214616 36604 418160 36632
rect 214616 36592 214622 36604
rect 418154 36592 418160 36604
rect 418212 36592 418218 36644
rect 236086 36524 236092 36576
rect 236144 36564 236150 36576
rect 506566 36564 506572 36576
rect 236144 36536 506572 36564
rect 236144 36524 236150 36536
rect 506566 36524 506572 36536
rect 506624 36524 506630 36576
rect 191190 35436 191196 35488
rect 191248 35476 191254 35488
rect 340874 35476 340880 35488
rect 191248 35448 340880 35476
rect 191248 35436 191254 35448
rect 340874 35436 340880 35448
rect 340932 35436 340938 35488
rect 183646 35368 183652 35420
rect 183704 35408 183710 35420
rect 338114 35408 338120 35420
rect 183704 35380 338120 35408
rect 183704 35368 183710 35380
rect 338114 35368 338120 35380
rect 338172 35368 338178 35420
rect 140958 35300 140964 35352
rect 141016 35340 141022 35352
rect 188430 35340 188436 35352
rect 141016 35312 188436 35340
rect 141016 35300 141022 35312
rect 188430 35300 188436 35312
rect 188488 35300 188494 35352
rect 254026 35300 254032 35352
rect 254084 35340 254090 35352
rect 564618 35340 564624 35352
rect 254084 35312 564624 35340
rect 254084 35300 254090 35312
rect 564618 35300 564624 35312
rect 564676 35300 564682 35352
rect 147858 35232 147864 35284
rect 147916 35272 147922 35284
rect 222378 35272 222384 35284
rect 147916 35244 222384 35272
rect 147916 35232 147922 35244
rect 222378 35232 222384 35244
rect 222436 35232 222442 35284
rect 256694 35232 256700 35284
rect 256752 35272 256758 35284
rect 572806 35272 572812 35284
rect 256752 35244 572812 35272
rect 256752 35232 256758 35244
rect 572806 35232 572812 35244
rect 572864 35232 572870 35284
rect 151906 35164 151912 35216
rect 151964 35204 151970 35216
rect 233418 35204 233424 35216
rect 151964 35176 233424 35204
rect 151964 35164 151970 35176
rect 233418 35164 233424 35176
rect 233476 35164 233482 35216
rect 256786 35164 256792 35216
rect 256844 35204 256850 35216
rect 575474 35204 575480 35216
rect 256844 35176 575480 35204
rect 256844 35164 256850 35176
rect 575474 35164 575480 35176
rect 575532 35164 575538 35216
rect 180978 34008 180984 34060
rect 181036 34048 181042 34060
rect 327074 34048 327080 34060
rect 181036 34020 327080 34048
rect 181036 34008 181042 34020
rect 327074 34008 327080 34020
rect 327132 34008 327138 34060
rect 182266 33940 182272 33992
rect 182324 33980 182330 33992
rect 331214 33980 331220 33992
rect 182324 33952 331220 33980
rect 182324 33940 182330 33952
rect 331214 33940 331220 33952
rect 331272 33940 331278 33992
rect 182358 33872 182364 33924
rect 182416 33912 182422 33924
rect 333974 33912 333980 33924
rect 182416 33884 333980 33912
rect 182416 33872 182422 33884
rect 333974 33872 333980 33884
rect 334032 33872 334038 33924
rect 213270 33804 213276 33856
rect 213328 33844 213334 33856
rect 415486 33844 415492 33856
rect 213328 33816 415492 33844
rect 213328 33804 213334 33816
rect 415486 33804 415492 33816
rect 415544 33804 415550 33856
rect 147766 33736 147772 33788
rect 147824 33776 147830 33788
rect 218238 33776 218244 33788
rect 147824 33748 218244 33776
rect 147824 33736 147830 33748
rect 218238 33736 218244 33748
rect 218296 33736 218302 33788
rect 226426 33736 226432 33788
rect 226484 33776 226490 33788
rect 477494 33776 477500 33788
rect 226484 33748 477500 33776
rect 226484 33736 226490 33748
rect 477494 33736 477500 33748
rect 477552 33736 477558 33788
rect 176838 32648 176844 32700
rect 176896 32688 176902 32700
rect 316034 32688 316040 32700
rect 176896 32660 316040 32688
rect 176896 32648 176902 32660
rect 316034 32648 316040 32660
rect 316092 32648 316098 32700
rect 178218 32580 178224 32632
rect 178276 32620 178282 32632
rect 320174 32620 320180 32632
rect 178276 32592 320180 32620
rect 178276 32580 178282 32592
rect 320174 32580 320180 32592
rect 320232 32580 320238 32632
rect 179506 32512 179512 32564
rect 179564 32552 179570 32564
rect 324406 32552 324412 32564
rect 179564 32524 324412 32552
rect 179564 32512 179570 32524
rect 324406 32512 324412 32524
rect 324464 32512 324470 32564
rect 213178 32444 213184 32496
rect 213236 32484 213242 32496
rect 411254 32484 411260 32496
rect 213236 32456 411260 32484
rect 213236 32444 213242 32456
rect 411254 32444 411260 32456
rect 411312 32444 411318 32496
rect 146478 32376 146484 32428
rect 146536 32416 146542 32428
rect 215294 32416 215300 32428
rect 146536 32388 215300 32416
rect 146536 32376 146542 32388
rect 215294 32376 215300 32388
rect 215352 32376 215358 32428
rect 218146 32376 218152 32428
rect 218204 32416 218210 32428
rect 448606 32416 448612 32428
rect 218204 32388 448612 32416
rect 218204 32376 218210 32388
rect 448606 32376 448612 32388
rect 448664 32376 448670 32428
rect 173986 31288 173992 31340
rect 174044 31328 174050 31340
rect 306374 31328 306380 31340
rect 174044 31300 306380 31328
rect 174044 31288 174050 31300
rect 306374 31288 306380 31300
rect 306432 31288 306438 31340
rect 175458 31220 175464 31272
rect 175516 31260 175522 31272
rect 309134 31260 309140 31272
rect 175516 31232 309140 31260
rect 175516 31220 175522 31232
rect 309134 31220 309140 31232
rect 309192 31220 309198 31272
rect 176746 31152 176752 31204
rect 176804 31192 176810 31204
rect 313274 31192 313280 31204
rect 176804 31164 313280 31192
rect 176804 31152 176810 31164
rect 313274 31152 313280 31164
rect 313332 31152 313338 31204
rect 139670 31084 139676 31136
rect 139728 31124 139734 31136
rect 174538 31124 174544 31136
rect 139728 31096 174544 31124
rect 139728 31084 139734 31096
rect 174538 31084 174544 31096
rect 174596 31084 174602 31136
rect 209130 31084 209136 31136
rect 209188 31124 209194 31136
rect 407114 31124 407120 31136
rect 209188 31096 407120 31124
rect 209188 31084 209194 31096
rect 407114 31084 407120 31096
rect 407172 31084 407178 31136
rect 143718 31016 143724 31068
rect 143776 31056 143782 31068
rect 208486 31056 208492 31068
rect 143776 31028 208492 31056
rect 143776 31016 143782 31028
rect 208486 31016 208492 31028
rect 208544 31016 208550 31068
rect 224954 31016 224960 31068
rect 225012 31056 225018 31068
rect 470594 31056 470600 31068
rect 225012 31028 470600 31056
rect 225012 31016 225018 31028
rect 470594 31016 470600 31028
rect 470652 31016 470658 31068
rect 165614 29928 165620 29980
rect 165672 29968 165678 29980
rect 277394 29968 277400 29980
rect 165672 29940 277400 29968
rect 165672 29928 165678 29940
rect 277394 29928 277400 29940
rect 277452 29928 277458 29980
rect 172790 29860 172796 29912
rect 172848 29900 172854 29912
rect 302234 29900 302240 29912
rect 172848 29872 302240 29900
rect 172848 29860 172854 29872
rect 302234 29860 302240 29872
rect 302292 29860 302298 29912
rect 195974 29792 195980 29844
rect 196032 29832 196038 29844
rect 375374 29832 375380 29844
rect 196032 29804 375380 29832
rect 196032 29792 196038 29804
rect 375374 29792 375380 29804
rect 375432 29792 375438 29844
rect 138198 29724 138204 29776
rect 138256 29764 138262 29776
rect 166350 29764 166356 29776
rect 138256 29736 166356 29764
rect 138256 29724 138262 29736
rect 166350 29724 166356 29736
rect 166408 29724 166414 29776
rect 251358 29724 251364 29776
rect 251416 29764 251422 29776
rect 557534 29764 557540 29776
rect 251416 29736 557540 29764
rect 251416 29724 251422 29736
rect 557534 29724 557540 29736
rect 557592 29724 557598 29776
rect 142430 29656 142436 29708
rect 142488 29696 142494 29708
rect 201586 29696 201592 29708
rect 142488 29668 201592 29696
rect 142488 29656 142494 29668
rect 201586 29656 201592 29668
rect 201644 29656 201650 29708
rect 252646 29656 252652 29708
rect 252704 29696 252710 29708
rect 561858 29696 561864 29708
rect 252704 29668 561864 29696
rect 252704 29656 252710 29668
rect 561858 29656 561864 29668
rect 561916 29656 561922 29708
rect 142338 29588 142344 29640
rect 142396 29628 142402 29640
rect 204254 29628 204260 29640
rect 142396 29600 204260 29628
rect 142396 29588 142402 29600
rect 204254 29588 204260 29600
rect 204312 29588 204318 29640
rect 255406 29588 255412 29640
rect 255464 29628 255470 29640
rect 568574 29628 568580 29640
rect 255464 29600 568580 29628
rect 255464 29588 255470 29600
rect 568574 29588 568580 29600
rect 568632 29588 568638 29640
rect 161566 28568 161572 28620
rect 161624 28608 161630 28620
rect 267826 28608 267832 28620
rect 161624 28580 267832 28608
rect 161624 28568 161630 28580
rect 267826 28568 267832 28580
rect 267884 28568 267890 28620
rect 164234 28500 164240 28552
rect 164292 28540 164298 28552
rect 274634 28540 274640 28552
rect 164292 28512 274640 28540
rect 164292 28500 164298 28512
rect 274634 28500 274640 28512
rect 274692 28500 274698 28552
rect 192570 28432 192576 28484
rect 192628 28472 192634 28484
rect 350534 28472 350540 28484
rect 192628 28444 350540 28472
rect 192628 28432 192634 28444
rect 350534 28432 350540 28444
rect 350592 28432 350598 28484
rect 244274 28364 244280 28416
rect 244332 28404 244338 28416
rect 532694 28404 532700 28416
rect 244332 28376 532700 28404
rect 244332 28364 244338 28376
rect 532694 28364 532700 28376
rect 532752 28364 532758 28416
rect 136910 28296 136916 28348
rect 136968 28336 136974 28348
rect 185026 28336 185032 28348
rect 136968 28308 185032 28336
rect 136968 28296 136974 28308
rect 185026 28296 185032 28308
rect 185084 28296 185090 28348
rect 249978 28296 249984 28348
rect 250036 28336 250042 28348
rect 550634 28336 550640 28348
rect 250036 28308 550640 28336
rect 250036 28296 250042 28308
rect 550634 28296 550640 28308
rect 550692 28296 550698 28348
rect 140866 28228 140872 28280
rect 140924 28268 140930 28280
rect 197446 28268 197452 28280
rect 140924 28240 197452 28268
rect 140924 28228 140930 28240
rect 197446 28228 197452 28240
rect 197504 28228 197510 28280
rect 251266 28228 251272 28280
rect 251324 28268 251330 28280
rect 554774 28268 554780 28280
rect 251324 28240 554780 28268
rect 251324 28228 251330 28240
rect 554774 28228 554780 28240
rect 554832 28228 554838 28280
rect 160094 27208 160100 27260
rect 160152 27248 160158 27260
rect 259638 27248 259644 27260
rect 160152 27220 259644 27248
rect 160152 27208 160158 27220
rect 259638 27208 259644 27220
rect 259696 27208 259702 27260
rect 161474 27140 161480 27192
rect 161532 27180 161538 27192
rect 263594 27180 263600 27192
rect 161532 27152 263600 27180
rect 161532 27140 161538 27152
rect 263594 27140 263600 27152
rect 263652 27140 263658 27192
rect 197354 27072 197360 27124
rect 197412 27112 197418 27124
rect 379514 27112 379520 27124
rect 197412 27084 379520 27112
rect 197412 27072 197418 27084
rect 379514 27072 379520 27084
rect 379572 27072 379578 27124
rect 132770 27004 132776 27056
rect 132828 27044 132834 27056
rect 160738 27044 160744 27056
rect 132828 27016 160744 27044
rect 132828 27004 132834 27016
rect 160738 27004 160744 27016
rect 160796 27004 160802 27056
rect 237374 27004 237380 27056
rect 237432 27044 237438 27056
rect 511994 27044 512000 27056
rect 237432 27016 512000 27044
rect 237432 27004 237438 27016
rect 511994 27004 512000 27016
rect 512052 27004 512058 27056
rect 139578 26936 139584 26988
rect 139636 26976 139642 26988
rect 193306 26976 193312 26988
rect 139636 26948 193312 26976
rect 139636 26936 139642 26948
rect 193306 26936 193312 26948
rect 193364 26936 193370 26988
rect 241606 26936 241612 26988
rect 241664 26976 241670 26988
rect 523126 26976 523132 26988
rect 241664 26948 523132 26976
rect 241664 26936 241670 26948
rect 523126 26936 523132 26948
rect 523184 26936 523190 26988
rect 150710 26868 150716 26920
rect 150768 26908 150774 26920
rect 229186 26908 229192 26920
rect 150768 26880 229192 26908
rect 150768 26868 150774 26880
rect 229186 26868 229192 26880
rect 229244 26868 229250 26920
rect 241698 26868 241704 26920
rect 241756 26908 241762 26920
rect 525794 26908 525800 26920
rect 241756 26880 525800 26908
rect 241756 26868 241762 26880
rect 525794 26868 525800 26880
rect 525852 26868 525858 26920
rect 156138 25848 156144 25900
rect 156196 25888 156202 25900
rect 249978 25888 249984 25900
rect 156196 25860 249984 25888
rect 156196 25848 156202 25860
rect 249978 25848 249984 25860
rect 250036 25848 250042 25900
rect 157426 25780 157432 25832
rect 157484 25820 157490 25832
rect 252646 25820 252652 25832
rect 157484 25792 252652 25820
rect 157484 25780 157490 25792
rect 252646 25780 252652 25792
rect 252704 25780 252710 25832
rect 186314 25712 186320 25764
rect 186372 25752 186378 25764
rect 343634 25752 343640 25764
rect 186372 25724 343640 25752
rect 186372 25712 186378 25724
rect 343634 25712 343640 25724
rect 343692 25712 343698 25764
rect 233326 25644 233332 25696
rect 233384 25684 233390 25696
rect 498286 25684 498292 25696
rect 233384 25656 498292 25684
rect 233384 25644 233390 25656
rect 498286 25644 498292 25656
rect 498344 25644 498350 25696
rect 234798 25576 234804 25628
rect 234856 25616 234862 25628
rect 500954 25616 500960 25628
rect 234856 25588 500960 25616
rect 234856 25576 234862 25588
rect 500954 25576 500960 25588
rect 501012 25576 501018 25628
rect 138106 25508 138112 25560
rect 138164 25548 138170 25560
rect 190638 25548 190644 25560
rect 138164 25520 190644 25548
rect 138164 25508 138170 25520
rect 190638 25508 190644 25520
rect 190696 25508 190702 25560
rect 235994 25508 236000 25560
rect 236052 25548 236058 25560
rect 507854 25548 507860 25560
rect 236052 25520 507860 25548
rect 236052 25508 236058 25520
rect 507854 25508 507860 25520
rect 507912 25508 507918 25560
rect 154758 24488 154764 24540
rect 154816 24528 154822 24540
rect 242986 24528 242992 24540
rect 154816 24500 242992 24528
rect 154816 24488 154822 24500
rect 242986 24488 242992 24500
rect 243044 24488 243050 24540
rect 156046 24420 156052 24472
rect 156104 24460 156110 24472
rect 245838 24460 245844 24472
rect 156104 24432 245844 24460
rect 156104 24420 156110 24432
rect 245838 24420 245844 24432
rect 245896 24420 245902 24472
rect 212534 24352 212540 24404
rect 212592 24392 212598 24404
rect 429194 24392 429200 24404
rect 212592 24364 429200 24392
rect 212592 24352 212598 24364
rect 429194 24352 429200 24364
rect 429252 24352 429258 24404
rect 230658 24284 230664 24336
rect 230716 24324 230722 24336
rect 487154 24324 487160 24336
rect 230716 24296 487160 24324
rect 230716 24284 230722 24296
rect 487154 24284 487160 24296
rect 487212 24284 487218 24336
rect 230750 24216 230756 24268
rect 230808 24256 230814 24268
rect 489914 24256 489920 24268
rect 230808 24228 489920 24256
rect 230808 24216 230814 24228
rect 489914 24216 489920 24228
rect 489972 24216 489978 24268
rect 134518 24148 134524 24200
rect 134576 24188 134582 24200
rect 166994 24188 167000 24200
rect 134576 24160 167000 24188
rect 134576 24148 134582 24160
rect 166994 24148 167000 24160
rect 167052 24148 167058 24200
rect 231946 24148 231952 24200
rect 232004 24188 232010 24200
rect 494054 24188 494060 24200
rect 232004 24160 494060 24188
rect 232004 24148 232010 24160
rect 494054 24148 494060 24160
rect 494112 24148 494118 24200
rect 136818 24080 136824 24132
rect 136876 24120 136882 24132
rect 183646 24120 183652 24132
rect 136876 24092 183652 24120
rect 136876 24080 136882 24092
rect 183646 24080 183652 24092
rect 183704 24080 183710 24132
rect 241514 24080 241520 24132
rect 241572 24120 241578 24132
rect 524414 24120 524420 24132
rect 241572 24092 524420 24120
rect 241572 24080 241578 24092
rect 524414 24080 524420 24092
rect 524472 24080 524478 24132
rect 110690 23400 110696 23452
rect 110748 23440 110754 23452
rect 113358 23440 113364 23452
rect 110748 23412 113364 23440
rect 110748 23400 110754 23412
rect 113358 23400 113364 23412
rect 113416 23400 113422 23452
rect 158806 22924 158812 22976
rect 158864 22964 158870 22976
rect 256694 22964 256700 22976
rect 158864 22936 256700 22964
rect 158864 22924 158870 22936
rect 256694 22924 256700 22936
rect 256752 22924 256758 22976
rect 218054 22856 218060 22908
rect 218112 22896 218118 22908
rect 449894 22896 449900 22908
rect 218112 22868 449900 22896
rect 218112 22856 218118 22868
rect 449894 22856 449900 22868
rect 449952 22856 449958 22908
rect 227806 22788 227812 22840
rect 227864 22828 227870 22840
rect 480254 22828 480260 22840
rect 227864 22800 480260 22828
rect 227864 22788 227870 22800
rect 480254 22788 480260 22800
rect 480312 22788 480318 22840
rect 53834 22720 53840 22772
rect 53892 22760 53898 22772
rect 96798 22760 96804 22772
rect 53892 22732 96804 22760
rect 53892 22720 53898 22732
rect 96798 22720 96804 22732
rect 96856 22720 96862 22772
rect 141418 22720 141424 22772
rect 141476 22760 141482 22772
rect 168466 22760 168472 22772
rect 141476 22732 168472 22760
rect 141476 22720 141482 22732
rect 168466 22720 168472 22732
rect 168524 22720 168530 22772
rect 240226 22720 240232 22772
rect 240284 22760 240290 22772
rect 521654 22760 521660 22772
rect 240284 22732 521660 22760
rect 240284 22720 240290 22732
rect 521654 22720 521660 22732
rect 521712 22720 521718 22772
rect 103882 22108 103888 22160
rect 103940 22148 103946 22160
rect 112070 22148 112076 22160
rect 103940 22120 112076 22148
rect 103940 22108 103946 22120
rect 112070 22108 112076 22120
rect 112128 22108 112134 22160
rect 178034 21632 178040 21684
rect 178092 21672 178098 21684
rect 318794 21672 318800 21684
rect 178092 21644 318800 21672
rect 178092 21632 178098 21644
rect 318794 21632 318800 21644
rect 318852 21632 318858 21684
rect 182174 21564 182180 21616
rect 182232 21604 182238 21616
rect 332686 21604 332692 21616
rect 182232 21576 332692 21604
rect 182232 21564 182238 21576
rect 332686 21564 332692 21576
rect 332744 21564 332750 21616
rect 144178 21496 144184 21548
rect 144236 21536 144242 21548
rect 179506 21536 179512 21548
rect 144236 21508 179512 21536
rect 144236 21496 144242 21508
rect 179506 21496 179512 21508
rect 179564 21496 179570 21548
rect 183554 21496 183560 21548
rect 183612 21536 183618 21548
rect 336734 21536 336740 21548
rect 183612 21508 336740 21536
rect 183612 21496 183618 21508
rect 336734 21496 336740 21508
rect 336792 21496 336798 21548
rect 132678 21428 132684 21480
rect 132736 21468 132742 21480
rect 172790 21468 172796 21480
rect 132736 21440 172796 21468
rect 132736 21428 132742 21440
rect 172790 21428 172796 21440
rect 172848 21428 172854 21480
rect 184934 21428 184940 21480
rect 184992 21468 184998 21480
rect 340966 21468 340972 21480
rect 184992 21440 340972 21468
rect 184992 21428 184998 21440
rect 340966 21428 340972 21440
rect 341024 21428 341030 21480
rect 77294 21360 77300 21412
rect 77352 21400 77358 21412
rect 103790 21400 103796 21412
rect 77352 21372 103796 21400
rect 77352 21360 77358 21372
rect 103790 21360 103796 21372
rect 103848 21360 103854 21412
rect 134058 21360 134064 21412
rect 134116 21400 134122 21412
rect 176746 21400 176752 21412
rect 134116 21372 176752 21400
rect 134116 21360 134122 21372
rect 176746 21360 176752 21372
rect 176804 21360 176810 21412
rect 210418 21360 210424 21412
rect 210476 21400 210482 21412
rect 404354 21400 404360 21412
rect 210476 21372 404360 21400
rect 210476 21360 210482 21372
rect 404354 21360 404360 21372
rect 404412 21360 404418 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 560110 20652 560116 20664
rect 3476 20624 560116 20652
rect 3476 20612 3482 20624
rect 560110 20612 560116 20624
rect 560168 20612 560174 20664
rect 560938 20612 560944 20664
rect 560996 20652 561002 20664
rect 579982 20652 579988 20664
rect 560996 20624 579988 20652
rect 560996 20612 561002 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 172698 20204 172704 20256
rect 172756 20244 172762 20256
rect 300854 20244 300860 20256
rect 172756 20216 300860 20244
rect 172756 20204 172762 20216
rect 300854 20204 300860 20216
rect 300912 20204 300918 20256
rect 173894 20136 173900 20188
rect 173952 20176 173958 20188
rect 304994 20176 305000 20188
rect 173952 20148 305000 20176
rect 173952 20136 173958 20148
rect 304994 20136 305000 20148
rect 305052 20136 305058 20188
rect 133966 20068 133972 20120
rect 134024 20108 134030 20120
rect 162118 20108 162124 20120
rect 134024 20080 162124 20108
rect 134024 20068 134030 20080
rect 162118 20068 162124 20080
rect 162176 20068 162182 20120
rect 175274 20068 175280 20120
rect 175332 20108 175338 20120
rect 307846 20108 307852 20120
rect 175332 20080 307852 20108
rect 175332 20068 175338 20080
rect 307846 20068 307852 20080
rect 307904 20068 307910 20120
rect 132586 20000 132592 20052
rect 132644 20040 132650 20052
rect 160830 20040 160836 20052
rect 132644 20012 160836 20040
rect 132644 20000 132650 20012
rect 160830 20000 160836 20012
rect 160888 20000 160894 20052
rect 175366 20000 175372 20052
rect 175424 20040 175430 20052
rect 311894 20040 311900 20052
rect 175424 20012 311900 20040
rect 175424 20000 175430 20012
rect 311894 20000 311900 20012
rect 311952 20000 311958 20052
rect 98270 19932 98276 19984
rect 98328 19972 98334 19984
rect 110598 19972 110604 19984
rect 98328 19944 110604 19972
rect 98328 19932 98334 19944
rect 110598 19932 110604 19944
rect 110656 19932 110662 19984
rect 130010 19932 130016 19984
rect 130068 19972 130074 19984
rect 161474 19972 161480 19984
rect 130068 19944 161480 19972
rect 130068 19932 130074 19944
rect 161474 19932 161480 19944
rect 161532 19932 161538 19984
rect 207658 19932 207664 19984
rect 207716 19972 207722 19984
rect 397454 19972 397460 19984
rect 207716 19944 397460 19972
rect 207716 19932 207722 19944
rect 397454 19932 397460 19944
rect 397512 19932 397518 19984
rect 179414 18844 179420 18896
rect 179472 18884 179478 18896
rect 322934 18884 322940 18896
rect 179472 18856 322940 18884
rect 179472 18844 179478 18856
rect 322934 18844 322940 18856
rect 322992 18844 322998 18896
rect 188338 18776 188344 18828
rect 188396 18816 188402 18828
rect 238754 18816 238760 18828
rect 188396 18788 238760 18816
rect 188396 18776 188402 18788
rect 238754 18776 238760 18788
rect 238812 18776 238818 18828
rect 245746 18776 245752 18828
rect 245804 18816 245810 18828
rect 539686 18816 539692 18828
rect 245804 18788 539692 18816
rect 245804 18776 245810 18788
rect 539686 18776 539692 18788
rect 539744 18776 539750 18828
rect 144914 18708 144920 18760
rect 144972 18748 144978 18760
rect 214006 18748 214012 18760
rect 144972 18720 214012 18748
rect 144972 18708 144978 18720
rect 214006 18708 214012 18720
rect 214064 18708 214070 18760
rect 252554 18708 252560 18760
rect 252612 18748 252618 18760
rect 560294 18748 560300 18760
rect 252612 18720 560300 18748
rect 252612 18708 252618 18720
rect 560294 18708 560300 18720
rect 560352 18708 560358 18760
rect 150618 18640 150624 18692
rect 150676 18680 150682 18692
rect 231946 18680 231952 18692
rect 150676 18652 231952 18680
rect 150676 18640 150682 18652
rect 231946 18640 231952 18652
rect 232004 18640 232010 18692
rect 255314 18640 255320 18692
rect 255372 18680 255378 18692
rect 567194 18680 567200 18692
rect 255372 18652 567200 18680
rect 255372 18640 255378 18652
rect 567194 18640 567200 18652
rect 567252 18640 567258 18692
rect 24854 18572 24860 18624
rect 24912 18612 24918 18624
rect 87138 18612 87144 18624
rect 24912 18584 87144 18612
rect 24912 18572 24918 18584
rect 87138 18572 87144 18584
rect 87196 18572 87202 18624
rect 124490 18572 124496 18624
rect 124548 18612 124554 18624
rect 144914 18612 144920 18624
rect 124548 18584 144920 18612
rect 124548 18572 124554 18584
rect 144914 18572 144920 18584
rect 144972 18572 144978 18624
rect 151814 18572 151820 18624
rect 151872 18612 151878 18624
rect 234798 18612 234804 18624
rect 151872 18584 234804 18612
rect 151872 18572 151878 18584
rect 234798 18572 234804 18584
rect 234856 18572 234862 18624
rect 258074 18572 258080 18624
rect 258132 18612 258138 18624
rect 578234 18612 578240 18624
rect 258132 18584 578240 18612
rect 258132 18572 258138 18584
rect 578234 18572 578240 18584
rect 578292 18572 578298 18624
rect 180886 17484 180892 17536
rect 180944 17524 180950 17536
rect 325694 17524 325700 17536
rect 180944 17496 325700 17524
rect 180944 17484 180950 17496
rect 325694 17484 325700 17496
rect 325752 17484 325758 17536
rect 60734 17416 60740 17468
rect 60792 17456 60798 17468
rect 98178 17456 98184 17468
rect 60792 17428 98184 17456
rect 60792 17416 60798 17428
rect 98178 17416 98184 17428
rect 98236 17416 98242 17468
rect 123018 17416 123024 17468
rect 123076 17456 123082 17468
rect 142338 17456 142344 17468
rect 123076 17428 142344 17456
rect 123076 17416 123082 17428
rect 142338 17416 142344 17428
rect 142396 17416 142402 17468
rect 231854 17416 231860 17468
rect 231912 17456 231918 17468
rect 492674 17456 492680 17468
rect 231912 17428 492680 17456
rect 231912 17416 231918 17428
rect 492674 17416 492680 17428
rect 492732 17416 492738 17468
rect 45554 17348 45560 17400
rect 45612 17388 45618 17400
rect 94038 17388 94044 17400
rect 45612 17360 94044 17388
rect 45612 17348 45618 17360
rect 94038 17348 94044 17360
rect 94096 17348 94102 17400
rect 139486 17348 139492 17400
rect 139544 17388 139550 17400
rect 195974 17388 195980 17400
rect 139544 17360 195980 17388
rect 139544 17348 139550 17360
rect 195974 17348 195980 17360
rect 196032 17348 196038 17400
rect 233234 17348 233240 17400
rect 233292 17388 233298 17400
rect 496814 17388 496820 17400
rect 233292 17360 496820 17388
rect 233292 17348 233298 17360
rect 496814 17348 496820 17360
rect 496872 17348 496878 17400
rect 38654 17280 38660 17332
rect 38712 17320 38718 17332
rect 91278 17320 91284 17332
rect 38712 17292 91284 17320
rect 38712 17280 38718 17292
rect 91278 17280 91284 17292
rect 91336 17280 91342 17332
rect 140774 17280 140780 17332
rect 140832 17320 140838 17332
rect 200206 17320 200212 17332
rect 140832 17292 200212 17320
rect 140832 17280 140838 17292
rect 200206 17280 200212 17292
rect 200264 17280 200270 17332
rect 234706 17280 234712 17332
rect 234764 17320 234770 17332
rect 499574 17320 499580 17332
rect 234764 17292 499580 17320
rect 234764 17280 234770 17292
rect 499574 17280 499580 17292
rect 499632 17280 499638 17332
rect 15194 17212 15200 17264
rect 15252 17252 15258 17264
rect 84286 17252 84292 17264
rect 15252 17224 84292 17252
rect 15252 17212 15258 17224
rect 84286 17212 84292 17224
rect 84344 17212 84350 17264
rect 142246 17212 142252 17264
rect 142304 17252 142310 17264
rect 202874 17252 202880 17264
rect 142304 17224 202880 17252
rect 142304 17212 142310 17224
rect 202874 17212 202880 17224
rect 202932 17212 202938 17264
rect 234614 17212 234620 17264
rect 234672 17252 234678 17264
rect 503714 17252 503720 17264
rect 234672 17224 503720 17252
rect 234672 17212 234678 17224
rect 503714 17212 503720 17224
rect 503772 17212 503778 17264
rect 191098 16124 191104 16176
rect 191156 16164 191162 16176
rect 348050 16164 348056 16176
rect 191156 16136 348056 16164
rect 191156 16124 191162 16136
rect 348050 16124 348056 16136
rect 348108 16124 348114 16176
rect 74994 16056 75000 16108
rect 75052 16096 75058 16108
rect 100018 16096 100024 16108
rect 75052 16068 100024 16096
rect 75052 16056 75058 16068
rect 100018 16056 100024 16068
rect 100076 16056 100082 16108
rect 166258 16056 166264 16108
rect 166316 16096 166322 16108
rect 182174 16096 182180 16108
rect 166316 16068 182180 16096
rect 166316 16056 166322 16068
rect 182174 16056 182180 16068
rect 182232 16056 182238 16108
rect 205726 16056 205732 16108
rect 205784 16096 205790 16108
rect 407206 16096 407212 16108
rect 205784 16068 407212 16096
rect 205784 16056 205790 16068
rect 407206 16056 407212 16068
rect 407264 16056 407270 16108
rect 67634 15988 67640 16040
rect 67692 16028 67698 16040
rect 100938 16028 100944 16040
rect 67692 16000 100944 16028
rect 67692 15988 67698 16000
rect 100938 15988 100944 16000
rect 100996 15988 101002 16040
rect 136726 15988 136732 16040
rect 136784 16028 136790 16040
rect 170398 16028 170404 16040
rect 136784 16000 170404 16028
rect 136784 15988 136790 16000
rect 170398 15988 170404 16000
rect 170456 15988 170462 16040
rect 205818 15988 205824 16040
rect 205876 16028 205882 16040
rect 410794 16028 410800 16040
rect 205876 16000 410800 16028
rect 205876 15988 205882 16000
rect 410794 15988 410800 16000
rect 410852 15988 410858 16040
rect 31938 15920 31944 15972
rect 31996 15960 32002 15972
rect 89898 15960 89904 15972
rect 31996 15932 89904 15960
rect 31996 15920 32002 15932
rect 89898 15920 89904 15932
rect 89956 15920 89962 15972
rect 133874 15920 133880 15972
rect 133932 15960 133938 15972
rect 175458 15960 175464 15972
rect 133932 15932 175464 15960
rect 133932 15920 133938 15932
rect 175458 15920 175464 15932
rect 175516 15920 175522 15972
rect 208394 15920 208400 15972
rect 208452 15960 208458 15972
rect 417418 15960 417424 15972
rect 208452 15932 417424 15960
rect 208452 15920 208458 15932
rect 417418 15920 417424 15932
rect 417476 15920 417482 15972
rect 24210 15852 24216 15904
rect 24268 15892 24274 15904
rect 87046 15892 87052 15904
rect 24268 15864 87052 15892
rect 24268 15852 24274 15864
rect 87046 15852 87052 15864
rect 87104 15852 87110 15904
rect 122926 15852 122932 15904
rect 122984 15892 122990 15904
rect 138842 15892 138848 15904
rect 122984 15864 138848 15892
rect 122984 15852 122990 15864
rect 138842 15852 138848 15864
rect 138900 15852 138906 15904
rect 139394 15852 139400 15904
rect 139452 15892 139458 15904
rect 193398 15892 193404 15904
rect 139452 15864 193404 15892
rect 139452 15852 139458 15864
rect 193398 15852 193404 15864
rect 193456 15852 193462 15904
rect 223574 15852 223580 15904
rect 223632 15892 223638 15904
rect 467466 15892 467472 15904
rect 223632 15864 467472 15892
rect 223632 15852 223638 15864
rect 467466 15852 467472 15864
rect 467524 15852 467530 15904
rect 190546 14696 190552 14748
rect 190604 14736 190610 14748
rect 361114 14736 361120 14748
rect 190604 14708 361120 14736
rect 190604 14696 190610 14708
rect 361114 14696 361120 14708
rect 361172 14696 361178 14748
rect 56778 14628 56784 14680
rect 56836 14668 56842 14680
rect 96706 14668 96712 14680
rect 56836 14640 96712 14668
rect 56836 14628 56842 14640
rect 96706 14628 96712 14640
rect 96764 14628 96770 14680
rect 191834 14628 191840 14680
rect 191892 14668 191898 14680
rect 364610 14668 364616 14680
rect 191892 14640 364616 14668
rect 191892 14628 191898 14640
rect 364610 14628 364616 14640
rect 364668 14628 364674 14680
rect 53006 14560 53012 14612
rect 53064 14600 53070 14612
rect 93118 14600 93124 14612
rect 53064 14572 93124 14600
rect 53064 14560 53070 14572
rect 93118 14560 93124 14572
rect 93176 14560 93182 14612
rect 129826 14560 129832 14612
rect 129884 14600 129890 14612
rect 160646 14600 160652 14612
rect 129884 14572 160652 14600
rect 129884 14560 129890 14572
rect 160646 14560 160652 14572
rect 160704 14560 160710 14612
rect 193214 14560 193220 14612
rect 193272 14600 193278 14612
rect 367738 14600 367744 14612
rect 193272 14572 367744 14600
rect 193272 14560 193278 14572
rect 367738 14560 367744 14572
rect 367796 14560 367802 14612
rect 14274 14492 14280 14544
rect 14332 14532 14338 14544
rect 84194 14532 84200 14544
rect 14332 14504 84200 14532
rect 14332 14492 14338 14504
rect 84194 14492 84200 14504
rect 84252 14492 84258 14544
rect 129918 14492 129924 14544
rect 129976 14532 129982 14544
rect 164418 14532 164424 14544
rect 129976 14504 164424 14532
rect 129976 14492 129982 14504
rect 164418 14492 164424 14504
rect 164476 14492 164482 14544
rect 200114 14492 200120 14544
rect 200172 14532 200178 14544
rect 390646 14532 390652 14544
rect 200172 14504 390652 14532
rect 200172 14492 200178 14504
rect 390646 14492 390652 14504
rect 390704 14492 390710 14544
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 82998 14464 83004 14476
rect 9732 14436 83004 14464
rect 9732 14424 9738 14436
rect 82998 14424 83004 14436
rect 83056 14424 83062 14476
rect 85758 14424 85764 14476
rect 85816 14464 85822 14476
rect 101398 14464 101404 14476
rect 85816 14436 101404 14464
rect 85816 14424 85822 14436
rect 101398 14424 101404 14436
rect 101456 14424 101462 14476
rect 132494 14424 132500 14476
rect 132552 14464 132558 14476
rect 171962 14464 171968 14476
rect 132552 14436 171968 14464
rect 132552 14424 132558 14436
rect 171962 14424 171968 14436
rect 172020 14424 172026 14476
rect 222286 14424 222292 14476
rect 222344 14464 222350 14476
rect 463970 14464 463976 14476
rect 222344 14436 463976 14464
rect 222344 14424 222350 14436
rect 463970 14424 463976 14436
rect 464028 14424 464034 14476
rect 157334 13404 157340 13456
rect 157392 13444 157398 13456
rect 251266 13444 251272 13456
rect 157392 13416 251272 13444
rect 157392 13404 157398 13416
rect 251266 13404 251272 13416
rect 251324 13404 251330 13456
rect 172606 13336 172612 13388
rect 172664 13376 172670 13388
rect 299474 13376 299480 13388
rect 172664 13348 299480 13376
rect 172664 13336 172670 13348
rect 299474 13336 299480 13348
rect 299532 13336 299538 13388
rect 69842 13268 69848 13320
rect 69900 13308 69906 13320
rect 100846 13308 100852 13320
rect 69900 13280 100852 13308
rect 69900 13268 69906 13280
rect 100846 13268 100852 13280
rect 100904 13268 100910 13320
rect 158714 13268 158720 13320
rect 158772 13308 158778 13320
rect 255866 13308 255872 13320
rect 158772 13280 255872 13308
rect 158772 13268 158778 13280
rect 255866 13268 255872 13280
rect 255924 13268 255930 13320
rect 255958 13268 255964 13320
rect 256016 13308 256022 13320
rect 454034 13308 454040 13320
rect 256016 13280 454040 13308
rect 256016 13268 256022 13280
rect 454034 13268 454040 13280
rect 454092 13268 454098 13320
rect 41874 13200 41880 13252
rect 41932 13240 41938 13252
rect 92658 13240 92664 13252
rect 41932 13212 92664 13240
rect 41932 13200 41938 13212
rect 92658 13200 92664 13212
rect 92716 13200 92722 13252
rect 128354 13200 128360 13252
rect 128412 13240 128418 13252
rect 157794 13240 157800 13252
rect 128412 13212 157800 13240
rect 128412 13200 128418 13212
rect 157794 13200 157800 13212
rect 157852 13200 157858 13252
rect 222194 13200 222200 13252
rect 222252 13240 222258 13252
rect 459922 13240 459928 13252
rect 222252 13212 459928 13240
rect 222252 13200 222258 13212
rect 459922 13200 459928 13212
rect 459980 13200 459986 13252
rect 34514 13132 34520 13184
rect 34572 13172 34578 13184
rect 89806 13172 89812 13184
rect 34572 13144 89812 13172
rect 34572 13132 34578 13144
rect 89806 13132 89812 13144
rect 89864 13132 89870 13184
rect 128446 13132 128452 13184
rect 128504 13172 128510 13184
rect 158898 13172 158904 13184
rect 128504 13144 158904 13172
rect 128504 13132 128510 13144
rect 158898 13132 158904 13144
rect 158956 13132 158962 13184
rect 226334 13132 226340 13184
rect 226392 13172 226398 13184
rect 474090 13172 474096 13184
rect 226392 13144 474096 13172
rect 226392 13132 226398 13144
rect 474090 13132 474096 13144
rect 474148 13132 474154 13184
rect 27706 13064 27712 13116
rect 27764 13104 27770 13116
rect 88426 13104 88432 13116
rect 27764 13076 88432 13104
rect 27764 13064 27770 13076
rect 88426 13064 88432 13076
rect 88484 13064 88490 13116
rect 118878 13064 118884 13116
rect 118936 13104 118942 13116
rect 128170 13104 128176 13116
rect 118936 13076 128176 13104
rect 118936 13064 118942 13076
rect 128170 13064 128176 13076
rect 128228 13064 128234 13116
rect 129734 13064 129740 13116
rect 129792 13104 129798 13116
rect 163682 13104 163688 13116
rect 129792 13076 163688 13104
rect 129792 13064 129798 13076
rect 163682 13064 163688 13076
rect 163740 13064 163746 13116
rect 249886 13064 249892 13116
rect 249944 13104 249950 13116
rect 550266 13104 550272 13116
rect 249944 13076 550272 13104
rect 249944 13064 249950 13076
rect 550266 13064 550272 13076
rect 550324 13064 550330 13116
rect 143534 12724 143540 12776
rect 143592 12764 143598 12776
rect 143718 12764 143724 12776
rect 143592 12736 143724 12764
rect 143592 12724 143598 12736
rect 143718 12724 143724 12736
rect 143776 12724 143782 12776
rect 234798 12724 234804 12776
rect 234856 12764 234862 12776
rect 235810 12764 235816 12776
rect 234856 12736 235816 12764
rect 234856 12724 234862 12736
rect 235810 12724 235816 12736
rect 235868 12724 235874 12776
rect 176654 11976 176660 12028
rect 176712 12016 176718 12028
rect 316218 12016 316224 12028
rect 176712 11988 316224 12016
rect 176712 11976 176718 11988
rect 316218 11976 316224 11988
rect 316276 11976 316282 12028
rect 61562 11908 61568 11960
rect 61620 11948 61626 11960
rect 98086 11948 98092 11960
rect 61620 11920 98092 11948
rect 61620 11908 61626 11920
rect 98086 11908 98092 11920
rect 98144 11908 98150 11960
rect 230566 11908 230572 11960
rect 230624 11948 230630 11960
rect 490006 11948 490012 11960
rect 230624 11920 490012 11948
rect 230624 11908 230630 11920
rect 490006 11908 490012 11920
rect 490064 11908 490070 11960
rect 63218 11840 63224 11892
rect 63276 11880 63282 11892
rect 99466 11880 99472 11892
rect 63276 11852 99472 11880
rect 63276 11840 63282 11852
rect 99466 11840 99472 11852
rect 99524 11840 99530 11892
rect 125778 11840 125784 11892
rect 125836 11880 125842 11892
rect 150618 11880 150624 11892
rect 125836 11852 150624 11880
rect 125836 11840 125842 11852
rect 150618 11840 150624 11852
rect 150676 11840 150682 11892
rect 154666 11840 154672 11892
rect 154724 11880 154730 11892
rect 241698 11880 241704 11892
rect 154724 11852 241704 11880
rect 154724 11840 154730 11852
rect 241698 11840 241704 11852
rect 241756 11840 241762 11892
rect 245194 11880 245200 11892
rect 241992 11852 245200 11880
rect 44266 11772 44272 11824
rect 44324 11812 44330 11824
rect 92566 11812 92572 11824
rect 44324 11784 92572 11812
rect 44324 11772 44330 11784
rect 92566 11772 92572 11784
rect 92624 11772 92630 11824
rect 127158 11772 127164 11824
rect 127216 11812 127222 11824
rect 153746 11812 153752 11824
rect 127216 11784 153752 11812
rect 127216 11772 127222 11784
rect 153746 11772 153752 11784
rect 153804 11772 153810 11824
rect 154574 11772 154580 11824
rect 154632 11812 154638 11824
rect 241992 11812 242020 11852
rect 245194 11840 245200 11852
rect 245252 11840 245258 11892
rect 248506 11840 248512 11892
rect 248564 11880 248570 11892
rect 548610 11880 548616 11892
rect 248564 11852 548616 11880
rect 248564 11840 248570 11852
rect 548610 11840 548616 11852
rect 548668 11840 548674 11892
rect 154632 11784 242020 11812
rect 154632 11772 154638 11784
rect 242894 11772 242900 11824
rect 242952 11812 242958 11824
rect 244090 11812 244096 11824
rect 242952 11784 244096 11812
rect 242952 11772 242958 11784
rect 244090 11772 244096 11784
rect 244148 11772 244154 11824
rect 249794 11772 249800 11824
rect 249852 11812 249858 11824
rect 552658 11812 552664 11824
rect 249852 11784 552664 11812
rect 249852 11772 249858 11784
rect 552658 11772 552664 11784
rect 552716 11772 552722 11824
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 85666 11744 85672 11756
rect 18012 11716 85672 11744
rect 18012 11704 18018 11716
rect 85666 11704 85672 11716
rect 85724 11704 85730 11756
rect 89162 11704 89168 11756
rect 89220 11744 89226 11756
rect 105538 11744 105544 11756
rect 89220 11716 105544 11744
rect 89220 11704 89226 11716
rect 105538 11704 105544 11716
rect 105596 11704 105602 11756
rect 125686 11704 125692 11756
rect 125744 11744 125750 11756
rect 151814 11744 151820 11756
rect 125744 11716 151820 11744
rect 125744 11704 125750 11716
rect 151814 11704 151820 11716
rect 151872 11704 151878 11756
rect 155954 11704 155960 11756
rect 156012 11744 156018 11756
rect 248506 11744 248512 11756
rect 156012 11716 248512 11744
rect 156012 11704 156018 11716
rect 248506 11704 248512 11716
rect 248564 11704 248570 11756
rect 251174 11704 251180 11756
rect 251232 11744 251238 11756
rect 556246 11744 556252 11756
rect 251232 11716 556252 11744
rect 251232 11704 251238 11716
rect 556246 11704 556252 11716
rect 556304 11704 556310 11756
rect 117406 10956 117412 11008
rect 117464 10996 117470 11008
rect 120626 10996 120632 11008
rect 117464 10968 120632 10996
rect 117464 10956 117470 10968
rect 120626 10956 120632 10968
rect 120684 10956 120690 11008
rect 150526 10616 150532 10668
rect 150584 10656 150590 10668
rect 231026 10656 231032 10668
rect 150584 10628 231032 10656
rect 150584 10616 150590 10628
rect 231026 10616 231032 10628
rect 231084 10616 231090 10668
rect 192478 10548 192484 10600
rect 192536 10588 192542 10600
rect 357526 10588 357532 10600
rect 192536 10560 357532 10588
rect 192536 10548 192542 10560
rect 357526 10548 357532 10560
rect 357584 10548 357590 10600
rect 56042 10480 56048 10532
rect 56100 10520 56106 10532
rect 96614 10520 96620 10532
rect 56100 10492 96620 10520
rect 56100 10480 56106 10492
rect 96614 10480 96620 10492
rect 96672 10480 96678 10532
rect 220814 10480 220820 10532
rect 220872 10520 220878 10532
rect 456886 10520 456892 10532
rect 220872 10492 456892 10520
rect 220872 10480 220878 10492
rect 456886 10480 456892 10492
rect 456944 10480 456950 10532
rect 40218 10412 40224 10464
rect 40276 10452 40282 10464
rect 92750 10452 92756 10464
rect 40276 10424 92756 10452
rect 40276 10412 40282 10424
rect 92750 10412 92756 10424
rect 92808 10412 92814 10464
rect 129090 10412 129096 10464
rect 129148 10452 129154 10464
rect 143534 10452 143540 10464
rect 129148 10424 143540 10452
rect 129148 10412 129154 10424
rect 143534 10412 143540 10424
rect 143592 10412 143598 10464
rect 227714 10412 227720 10464
rect 227772 10452 227778 10464
rect 481726 10452 481732 10464
rect 227772 10424 481732 10452
rect 227772 10412 227778 10424
rect 481726 10412 481732 10424
rect 481784 10412 481790 10464
rect 13538 10344 13544 10396
rect 13596 10384 13602 10396
rect 82906 10384 82912 10396
rect 13596 10356 82912 10384
rect 13596 10344 13602 10356
rect 82906 10344 82912 10356
rect 82964 10344 82970 10396
rect 92566 10344 92572 10396
rect 92624 10384 92630 10396
rect 107010 10384 107016 10396
rect 92624 10356 107016 10384
rect 92624 10344 92630 10356
rect 107010 10344 107016 10356
rect 107068 10344 107074 10396
rect 122834 10344 122840 10396
rect 122892 10384 122898 10396
rect 141234 10384 141240 10396
rect 122892 10356 141240 10384
rect 122892 10344 122898 10356
rect 141234 10344 141240 10356
rect 141292 10344 141298 10396
rect 146386 10344 146392 10396
rect 146444 10384 146450 10396
rect 216858 10384 216864 10396
rect 146444 10356 216864 10384
rect 146444 10344 146450 10356
rect 216858 10344 216864 10356
rect 216916 10344 216922 10396
rect 229094 10344 229100 10396
rect 229152 10384 229158 10396
rect 484762 10384 484768 10396
rect 229152 10356 484768 10384
rect 229152 10344 229158 10356
rect 484762 10344 484768 10356
rect 484820 10344 484826 10396
rect 3602 10276 3608 10328
rect 3660 10316 3666 10328
rect 80146 10316 80152 10328
rect 3660 10288 80152 10316
rect 3660 10276 3666 10288
rect 80146 10276 80152 10288
rect 80204 10276 80210 10328
rect 87506 10276 87512 10328
rect 87564 10316 87570 10328
rect 106366 10316 106372 10328
rect 87564 10288 106372 10316
rect 87564 10276 87570 10288
rect 106366 10276 106372 10288
rect 106424 10276 106430 10328
rect 125594 10276 125600 10328
rect 125652 10316 125658 10328
rect 147858 10316 147864 10328
rect 125652 10288 147864 10316
rect 125652 10276 125658 10288
rect 147858 10276 147864 10288
rect 147916 10276 147922 10328
rect 149054 10276 149060 10328
rect 149112 10316 149118 10328
rect 227530 10316 227536 10328
rect 149112 10288 227536 10316
rect 149112 10276 149118 10288
rect 227530 10276 227536 10288
rect 227588 10276 227594 10328
rect 230474 10276 230480 10328
rect 230532 10316 230538 10328
rect 488810 10316 488816 10328
rect 230532 10288 488816 10316
rect 230532 10276 230538 10288
rect 488810 10276 488816 10288
rect 488868 10276 488874 10328
rect 116210 9596 116216 9648
rect 116268 9636 116274 9648
rect 118786 9636 118792 9648
rect 116268 9608 118792 9636
rect 116268 9596 116274 9608
rect 118786 9596 118792 9608
rect 118844 9596 118850 9648
rect 143626 9256 143632 9308
rect 143684 9296 143690 9308
rect 209774 9296 209780 9308
rect 143684 9268 209780 9296
rect 143684 9256 143690 9268
rect 209774 9256 209780 9268
rect 209832 9256 209838 9308
rect 86862 9188 86868 9240
rect 86920 9228 86926 9240
rect 106458 9228 106464 9240
rect 86920 9200 106464 9228
rect 86920 9188 86926 9200
rect 106458 9188 106464 9200
rect 106516 9188 106522 9240
rect 198734 9188 198740 9240
rect 198792 9228 198798 9240
rect 387150 9228 387156 9240
rect 198792 9200 387156 9228
rect 198792 9188 198798 9200
rect 387150 9188 387156 9200
rect 387208 9188 387214 9240
rect 72602 9120 72608 9172
rect 72660 9160 72666 9172
rect 102226 9160 102232 9172
rect 72660 9132 102232 9160
rect 72660 9120 72666 9132
rect 102226 9120 102232 9132
rect 102284 9120 102290 9172
rect 118878 9120 118884 9172
rect 118936 9160 118942 9172
rect 129366 9160 129372 9172
rect 118936 9132 129372 9160
rect 118936 9120 118942 9132
rect 129366 9120 129372 9132
rect 129424 9120 129430 9172
rect 201494 9120 201500 9172
rect 201552 9160 201558 9172
rect 395338 9160 395344 9172
rect 201552 9132 395344 9160
rect 201552 9120 201558 9132
rect 395338 9120 395344 9132
rect 395396 9120 395402 9172
rect 58434 9052 58440 9104
rect 58492 9092 58498 9104
rect 97994 9092 98000 9104
rect 58492 9064 98000 9092
rect 58492 9052 58498 9064
rect 97994 9052 98000 9064
rect 98052 9052 98058 9104
rect 124398 9052 124404 9104
rect 124456 9092 124462 9104
rect 144730 9092 144736 9104
rect 124456 9064 144736 9092
rect 124456 9052 124462 9064
rect 144730 9052 144736 9064
rect 144788 9052 144794 9104
rect 205634 9052 205640 9104
rect 205692 9092 205698 9104
rect 409598 9092 409604 9104
rect 205692 9064 409604 9092
rect 205692 9052 205698 9064
rect 409598 9052 409604 9064
rect 409656 9052 409662 9104
rect 30098 8984 30104 9036
rect 30156 9024 30162 9036
rect 88610 9024 88616 9036
rect 30156 8996 88616 9024
rect 30156 8984 30162 8996
rect 88610 8984 88616 8996
rect 88668 8984 88674 9036
rect 123478 8984 123484 9036
rect 123536 9024 123542 9036
rect 134150 9024 134156 9036
rect 123536 8996 134156 9024
rect 123536 8984 123542 8996
rect 134150 8984 134156 8996
rect 134208 8984 134214 9036
rect 142154 8984 142160 9036
rect 142212 9024 142218 9036
rect 202690 9024 202696 9036
rect 142212 8996 202696 9024
rect 142212 8984 142218 8996
rect 202690 8984 202696 8996
rect 202748 8984 202754 9036
rect 209866 8984 209872 9036
rect 209924 9024 209930 9036
rect 423766 9024 423772 9036
rect 209924 8996 423772 9024
rect 209924 8984 209930 8996
rect 423766 8984 423772 8996
rect 423824 8984 423830 9036
rect 26510 8916 26516 8968
rect 26568 8956 26574 8968
rect 86954 8956 86960 8968
rect 26568 8928 86960 8956
rect 26568 8916 26574 8928
rect 86954 8916 86960 8928
rect 87012 8916 87018 8968
rect 101030 8916 101036 8968
rect 101088 8956 101094 8968
rect 110506 8956 110512 8968
rect 101088 8928 110512 8956
rect 101088 8916 101094 8928
rect 110506 8916 110512 8928
rect 110564 8916 110570 8968
rect 122098 8916 122104 8968
rect 122156 8956 122162 8968
rect 132954 8956 132960 8968
rect 122156 8928 132960 8956
rect 122156 8916 122162 8928
rect 132954 8916 132960 8928
rect 133012 8916 133018 8968
rect 143718 8916 143724 8968
rect 143776 8956 143782 8968
rect 206186 8956 206192 8968
rect 143776 8928 206192 8956
rect 143776 8916 143782 8928
rect 206186 8916 206192 8928
rect 206244 8916 206250 8968
rect 219434 8916 219440 8968
rect 219492 8956 219498 8968
rect 453298 8956 453304 8968
rect 219492 8928 453304 8956
rect 219492 8916 219498 8928
rect 453298 8916 453304 8928
rect 453356 8916 453362 8968
rect 117314 8236 117320 8288
rect 117372 8276 117378 8288
rect 122282 8276 122288 8288
rect 117372 8248 122288 8276
rect 117372 8236 117378 8248
rect 122282 8236 122288 8248
rect 122340 8236 122346 8288
rect 82078 7828 82084 7880
rect 82136 7868 82142 7880
rect 97258 7868 97264 7880
rect 82136 7840 97264 7868
rect 82136 7828 82142 7840
rect 97258 7828 97264 7840
rect 97316 7828 97322 7880
rect 187694 7828 187700 7880
rect 187752 7868 187758 7880
rect 349246 7868 349252 7880
rect 187752 7840 349252 7868
rect 187752 7828 187758 7840
rect 349246 7828 349252 7840
rect 349304 7828 349310 7880
rect 47854 7760 47860 7812
rect 47912 7800 47918 7812
rect 93946 7800 93952 7812
rect 47912 7772 93952 7800
rect 47912 7760 47918 7772
rect 93946 7760 93952 7772
rect 94004 7760 94010 7812
rect 121546 7760 121552 7812
rect 121604 7800 121610 7812
rect 137646 7800 137652 7812
rect 121604 7772 137652 7800
rect 121604 7760 121610 7772
rect 137646 7760 137652 7772
rect 137704 7760 137710 7812
rect 187786 7760 187792 7812
rect 187844 7800 187850 7812
rect 352834 7800 352840 7812
rect 187844 7772 352840 7800
rect 187844 7760 187850 7772
rect 352834 7760 352840 7772
rect 352892 7760 352898 7812
rect 21818 7692 21824 7744
rect 21876 7732 21882 7744
rect 85850 7732 85856 7744
rect 21876 7704 85856 7732
rect 21876 7692 21882 7704
rect 85850 7692 85856 7704
rect 85908 7692 85914 7744
rect 97442 7692 97448 7744
rect 97500 7732 97506 7744
rect 109218 7732 109224 7744
rect 97500 7704 109224 7732
rect 97500 7692 97506 7704
rect 109218 7692 109224 7704
rect 109276 7692 109282 7744
rect 138014 7692 138020 7744
rect 138072 7732 138078 7744
rect 188522 7732 188528 7744
rect 138072 7704 188528 7732
rect 138072 7692 138078 7704
rect 188522 7692 188528 7704
rect 188580 7692 188586 7744
rect 190454 7692 190460 7744
rect 190512 7732 190518 7744
rect 359918 7732 359924 7744
rect 190512 7704 359924 7732
rect 190512 7692 190518 7704
rect 359918 7692 359924 7704
rect 359976 7692 359982 7744
rect 7650 7624 7656 7676
rect 7708 7664 7714 7676
rect 81618 7664 81624 7676
rect 7708 7636 81624 7664
rect 7708 7624 7714 7636
rect 81618 7624 81624 7636
rect 81676 7624 81682 7676
rect 90358 7624 90364 7676
rect 90416 7664 90422 7676
rect 107838 7664 107844 7676
rect 90416 7636 107844 7664
rect 90416 7624 90422 7636
rect 107838 7624 107844 7636
rect 107896 7624 107902 7676
rect 121638 7624 121644 7676
rect 121696 7664 121702 7676
rect 135254 7664 135260 7676
rect 121696 7636 135260 7664
rect 121696 7624 121702 7636
rect 135254 7624 135260 7636
rect 135312 7624 135318 7676
rect 136634 7624 136640 7676
rect 136692 7664 136698 7676
rect 187326 7664 187332 7676
rect 136692 7636 187332 7664
rect 136692 7624 136698 7636
rect 187326 7624 187332 7636
rect 187384 7624 187390 7676
rect 209038 7624 209044 7676
rect 209096 7664 209102 7676
rect 394234 7664 394240 7676
rect 209096 7636 394240 7664
rect 209096 7624 209102 7636
rect 394234 7624 394240 7636
rect 394292 7624 394298 7676
rect 2866 7556 2872 7608
rect 2924 7596 2930 7608
rect 80054 7596 80060 7608
rect 2924 7568 80060 7596
rect 2924 7556 2930 7568
rect 80054 7556 80060 7568
rect 80112 7556 80118 7608
rect 80882 7556 80888 7608
rect 80940 7596 80946 7608
rect 105078 7596 105084 7608
rect 80940 7568 105084 7596
rect 80940 7556 80946 7568
rect 105078 7556 105084 7568
rect 105136 7556 105142 7608
rect 130562 7556 130568 7608
rect 130620 7596 130626 7608
rect 561674 7596 561680 7608
rect 130620 7568 561680 7596
rect 130620 7556 130626 7568
rect 561674 7556 561680 7568
rect 561732 7556 561738 7608
rect 561306 6808 561312 6860
rect 561364 6848 561370 6860
rect 580166 6848 580172 6860
rect 561364 6820 580172 6848
rect 561364 6808 561370 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 169754 6400 169760 6452
rect 169812 6440 169818 6452
rect 292574 6440 292580 6452
rect 169812 6412 292580 6440
rect 169812 6400 169818 6412
rect 292574 6400 292580 6412
rect 292632 6400 292638 6452
rect 77386 6332 77392 6384
rect 77444 6372 77450 6384
rect 103698 6372 103704 6384
rect 77444 6344 103704 6372
rect 77444 6332 77450 6344
rect 103698 6332 103704 6344
rect 103756 6332 103762 6384
rect 131206 6332 131212 6384
rect 131264 6372 131270 6384
rect 169570 6372 169576 6384
rect 131264 6344 169576 6372
rect 131264 6332 131270 6344
rect 169570 6332 169576 6344
rect 169628 6332 169634 6384
rect 172514 6332 172520 6384
rect 172572 6372 172578 6384
rect 299658 6372 299664 6384
rect 172572 6344 299664 6372
rect 172572 6332 172578 6344
rect 299658 6332 299664 6344
rect 299716 6332 299722 6384
rect 48958 6264 48964 6316
rect 49016 6304 49022 6316
rect 93854 6304 93860 6316
rect 49016 6276 93860 6304
rect 49016 6264 49022 6276
rect 93854 6264 93860 6276
rect 93912 6264 93918 6316
rect 126974 6264 126980 6316
rect 127032 6304 127038 6316
rect 127158 6304 127164 6316
rect 127032 6276 127164 6304
rect 127032 6264 127038 6276
rect 127158 6264 127164 6276
rect 127216 6264 127222 6316
rect 203518 6264 203524 6316
rect 203576 6304 203582 6316
rect 383562 6304 383568 6316
rect 203576 6276 383568 6304
rect 203576 6264 203582 6276
rect 383562 6264 383568 6276
rect 383620 6264 383626 6316
rect 33594 6196 33600 6248
rect 33652 6236 33658 6248
rect 89714 6236 89720 6248
rect 33652 6208 89720 6236
rect 33652 6196 33658 6208
rect 89714 6196 89720 6208
rect 89772 6196 89778 6248
rect 91554 6196 91560 6248
rect 91612 6236 91618 6248
rect 107746 6236 107752 6248
rect 91612 6208 107752 6236
rect 91612 6196 91618 6208
rect 107746 6196 107752 6208
rect 107804 6196 107810 6248
rect 131114 6196 131120 6248
rect 131172 6236 131178 6248
rect 166074 6236 166080 6248
rect 131172 6208 166080 6236
rect 131172 6196 131178 6208
rect 166074 6196 166080 6208
rect 166132 6196 166138 6248
rect 168374 6196 168380 6248
rect 168432 6236 168438 6248
rect 288986 6236 288992 6248
rect 168432 6208 288992 6236
rect 168432 6196 168438 6208
rect 288986 6196 288992 6208
rect 289044 6196 289050 6248
rect 289078 6196 289084 6248
rect 289136 6236 289142 6248
rect 475746 6236 475752 6248
rect 289136 6208 475752 6236
rect 289136 6196 289142 6208
rect 475746 6196 475752 6208
rect 475804 6196 475810 6248
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 81526 6168 81532 6180
rect 8812 6140 81532 6168
rect 8812 6128 8818 6140
rect 81526 6128 81532 6140
rect 81584 6128 81590 6180
rect 84470 6128 84476 6180
rect 84528 6168 84534 6180
rect 104986 6168 104992 6180
rect 84528 6140 104992 6168
rect 84528 6128 84534 6140
rect 104986 6128 104992 6140
rect 105044 6128 105050 6180
rect 126974 6128 126980 6180
rect 127032 6168 127038 6180
rect 561766 6168 561772 6180
rect 127032 6140 561772 6168
rect 127032 6128 127038 6140
rect 561766 6128 561772 6140
rect 561824 6128 561830 6180
rect 127066 5924 127072 5976
rect 127124 5964 127130 5976
rect 128354 5964 128360 5976
rect 127124 5936 128360 5964
rect 127124 5924 127130 5936
rect 128354 5924 128360 5936
rect 128412 5924 128418 5976
rect 126238 5516 126244 5568
rect 126296 5556 126302 5568
rect 131758 5556 131764 5568
rect 126296 5528 131764 5556
rect 126296 5516 126302 5528
rect 131758 5516 131764 5528
rect 131816 5516 131822 5568
rect 83274 5108 83280 5160
rect 83332 5148 83338 5160
rect 105170 5148 105176 5160
rect 83332 5120 105176 5148
rect 83332 5108 83338 5120
rect 105170 5108 105176 5120
rect 105228 5108 105234 5160
rect 187050 5108 187056 5160
rect 187108 5148 187114 5160
rect 225138 5148 225144 5160
rect 187108 5120 225144 5148
rect 187108 5108 187114 5120
rect 225138 5108 225144 5120
rect 225196 5108 225202 5160
rect 79686 5040 79692 5092
rect 79744 5080 79750 5092
rect 103606 5080 103612 5092
rect 79744 5052 103612 5080
rect 79744 5040 79750 5052
rect 103606 5040 103612 5052
rect 103664 5040 103670 5092
rect 180794 5040 180800 5092
rect 180852 5080 180858 5092
rect 330386 5080 330392 5092
rect 180852 5052 330392 5080
rect 180852 5040 180858 5052
rect 330386 5040 330392 5052
rect 330444 5040 330450 5092
rect 76190 4972 76196 5024
rect 76248 5012 76254 5024
rect 103514 5012 103520 5024
rect 76248 4984 103520 5012
rect 76248 4972 76254 4984
rect 103514 4972 103520 4984
rect 103572 4972 103578 5024
rect 213914 4972 213920 5024
rect 213972 5012 213978 5024
rect 437934 5012 437940 5024
rect 213972 4984 437940 5012
rect 213972 4972 213978 4984
rect 437934 4972 437940 4984
rect 437992 4972 437998 5024
rect 519538 5012 519544 5024
rect 509206 4984 519544 5012
rect 69106 4904 69112 4956
rect 69164 4944 69170 4956
rect 100938 4944 100944 4956
rect 69164 4916 100944 4944
rect 69164 4904 69170 4916
rect 100938 4904 100944 4916
rect 100996 4904 101002 4956
rect 118694 4904 118700 4956
rect 118752 4944 118758 4956
rect 125870 4944 125876 4956
rect 118752 4916 125876 4944
rect 118752 4904 118758 4916
rect 125870 4904 125876 4916
rect 125928 4904 125934 4956
rect 128998 4904 129004 4956
rect 129056 4944 129062 4956
rect 140038 4944 140044 4956
rect 129056 4916 140044 4944
rect 129056 4904 129062 4916
rect 140038 4904 140044 4916
rect 140096 4904 140102 4956
rect 146294 4904 146300 4956
rect 146352 4944 146358 4956
rect 218054 4944 218060 4956
rect 146352 4916 218060 4944
rect 146352 4904 146358 4916
rect 218054 4904 218060 4916
rect 218112 4904 218118 4956
rect 240134 4904 240140 4956
rect 240192 4944 240198 4956
rect 509206 4944 509234 4984
rect 519538 4972 519544 4984
rect 519596 4972 519602 5024
rect 240192 4916 509234 4944
rect 240192 4904 240198 4916
rect 65610 4836 65616 4888
rect 65668 4876 65674 4888
rect 99650 4876 99656 4888
rect 65668 4848 99656 4876
rect 65668 4836 65674 4848
rect 99650 4836 99656 4848
rect 99708 4836 99714 4888
rect 121454 4836 121460 4888
rect 121512 4876 121518 4888
rect 136450 4876 136456 4888
rect 121512 4848 136456 4876
rect 121512 4836 121518 4848
rect 136450 4836 136456 4848
rect 136508 4836 136514 4888
rect 147674 4836 147680 4888
rect 147732 4876 147738 4888
rect 221550 4876 221556 4888
rect 147732 4848 221556 4876
rect 147732 4836 147738 4848
rect 221550 4836 221556 4848
rect 221608 4836 221614 4888
rect 245654 4836 245660 4888
rect 245712 4876 245718 4888
rect 537202 4876 537208 4888
rect 245712 4848 537208 4876
rect 245712 4836 245718 4848
rect 537202 4836 537208 4848
rect 537260 4836 537266 4888
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 83090 4808 83096 4820
rect 12400 4780 83096 4808
rect 12400 4768 12406 4780
rect 83090 4768 83096 4780
rect 83148 4768 83154 4820
rect 124306 4768 124312 4820
rect 124364 4808 124370 4820
rect 147122 4808 147128 4820
rect 124364 4780 147128 4808
rect 124364 4768 124370 4780
rect 147122 4768 147128 4780
rect 147180 4768 147186 4820
rect 150434 4768 150440 4820
rect 150492 4808 150498 4820
rect 228726 4808 228732 4820
rect 150492 4780 228732 4808
rect 150492 4768 150498 4780
rect 228726 4768 228732 4780
rect 228784 4768 228790 4820
rect 248414 4768 248420 4820
rect 248472 4808 248478 4820
rect 547874 4808 547880 4820
rect 248472 4780 547880 4808
rect 248472 4768 248478 4780
rect 547874 4768 547880 4780
rect 547932 4768 547938 4820
rect 105722 4156 105728 4208
rect 105780 4196 105786 4208
rect 111978 4196 111984 4208
rect 105780 4168 111984 4196
rect 105780 4156 105786 4168
rect 111978 4156 111984 4168
rect 112036 4156 112042 4208
rect 64322 4088 64328 4140
rect 64380 4128 64386 4140
rect 65518 4128 65524 4140
rect 64380 4100 65524 4128
rect 64380 4088 64386 4100
rect 65518 4088 65524 4100
rect 65576 4088 65582 4140
rect 119338 4088 119344 4140
rect 119396 4128 119402 4140
rect 123478 4128 123484 4140
rect 119396 4100 123484 4128
rect 119396 4088 119402 4100
rect 123478 4088 123484 4100
rect 123536 4088 123542 4140
rect 170398 3748 170404 3800
rect 170456 3788 170462 3800
rect 170456 3760 171134 3788
rect 170456 3748 170462 3760
rect 162118 3680 162124 3732
rect 162176 3720 162182 3732
rect 162176 3692 170996 3720
rect 162176 3680 162182 3692
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 28258 3652 28264 3664
rect 20680 3624 28264 3652
rect 20680 3612 20686 3624
rect 28258 3612 28264 3624
rect 28316 3612 28322 3664
rect 109678 3652 109684 3664
rect 103486 3624 109684 3652
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 15838 3584 15844 3596
rect 11204 3556 15844 3584
rect 11204 3544 11210 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 43070 3544 43076 3596
rect 43128 3584 43134 3596
rect 53098 3584 53104 3596
rect 43128 3556 53104 3584
rect 43128 3544 43134 3556
rect 53098 3544 53104 3556
rect 53156 3544 53162 3596
rect 99834 3544 99840 3596
rect 99892 3584 99898 3596
rect 103486 3584 103514 3624
rect 109678 3612 109684 3624
rect 109736 3612 109742 3664
rect 160738 3612 160744 3664
rect 160796 3652 160802 3664
rect 160796 3624 161474 3652
rect 160796 3612 160802 3624
rect 108298 3584 108304 3596
rect 99892 3556 103514 3584
rect 104176 3556 108304 3584
rect 99892 3544 99898 3556
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 10318 3516 10324 3528
rect 5316 3488 10324 3516
rect 5316 3476 5322 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 28902 3476 28908 3528
rect 28960 3516 28966 3528
rect 32398 3516 32404 3528
rect 28960 3488 32404 3516
rect 28960 3476 28966 3488
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 44174 3476 44180 3528
rect 44232 3516 44238 3528
rect 45094 3516 45100 3528
rect 44232 3488 45100 3516
rect 44232 3476 44238 3488
rect 45094 3476 45100 3488
rect 45152 3476 45158 3528
rect 50338 3516 50344 3528
rect 45296 3488 50344 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 6512 3420 26234 3448
rect 6512 3408 6518 3420
rect 26206 3312 26234 3420
rect 35986 3340 35992 3392
rect 36044 3380 36050 3392
rect 45296 3380 45324 3488
rect 50338 3476 50344 3488
rect 50396 3476 50402 3528
rect 102134 3476 102140 3528
rect 102192 3516 102198 3528
rect 103330 3516 103336 3528
rect 102192 3488 103336 3516
rect 102192 3476 102198 3488
rect 103330 3476 103336 3488
rect 103388 3476 103394 3528
rect 103422 3476 103428 3528
rect 103480 3516 103486 3528
rect 104176 3516 104204 3556
rect 108298 3544 108304 3556
rect 108356 3544 108362 3596
rect 109310 3544 109316 3596
rect 109368 3584 109374 3596
rect 111058 3584 111064 3596
rect 109368 3556 111064 3584
rect 109368 3544 109374 3556
rect 111058 3544 111064 3556
rect 111116 3544 111122 3596
rect 128354 3544 128360 3596
rect 128412 3584 128418 3596
rect 153010 3584 153016 3596
rect 128412 3556 153016 3584
rect 128412 3544 128418 3556
rect 153010 3544 153016 3556
rect 153068 3544 153074 3596
rect 160830 3544 160836 3596
rect 160888 3544 160894 3596
rect 161446 3584 161474 3624
rect 170766 3584 170772 3596
rect 161446 3556 170772 3584
rect 170766 3544 170772 3556
rect 170824 3544 170830 3596
rect 170968 3584 170996 3692
rect 171106 3652 171134 3760
rect 407758 3748 407764 3800
rect 407816 3788 407822 3800
rect 461578 3788 461584 3800
rect 407816 3760 461584 3788
rect 407816 3748 407822 3760
rect 461578 3748 461584 3760
rect 461636 3748 461642 3800
rect 188430 3680 188436 3732
rect 188488 3720 188494 3732
rect 199102 3720 199108 3732
rect 188488 3692 199108 3720
rect 188488 3680 188494 3692
rect 199102 3680 199108 3692
rect 199160 3680 199166 3732
rect 411990 3680 411996 3732
rect 412048 3720 412054 3732
rect 468662 3720 468668 3732
rect 412048 3692 468668 3720
rect 412048 3680 412054 3692
rect 468662 3680 468668 3692
rect 468720 3680 468726 3732
rect 186130 3652 186136 3664
rect 171106 3624 186136 3652
rect 186130 3612 186136 3624
rect 186188 3612 186194 3664
rect 193306 3612 193312 3664
rect 193364 3652 193370 3664
rect 194410 3652 194416 3664
rect 193364 3624 194416 3652
rect 193364 3612 193370 3624
rect 194410 3612 194416 3624
rect 194468 3612 194474 3664
rect 258718 3612 258724 3664
rect 258776 3652 258782 3664
rect 258776 3624 259592 3652
rect 258776 3612 258782 3624
rect 177850 3584 177856 3596
rect 170968 3556 177856 3584
rect 177850 3544 177856 3556
rect 177908 3544 177914 3596
rect 186958 3544 186964 3596
rect 187016 3584 187022 3596
rect 207382 3584 207388 3596
rect 187016 3556 207388 3584
rect 187016 3544 187022 3556
rect 207382 3544 207388 3556
rect 207440 3544 207446 3596
rect 210510 3544 210516 3596
rect 210568 3584 210574 3596
rect 212166 3584 212172 3596
rect 210568 3556 212172 3584
rect 210568 3544 210574 3556
rect 212166 3544 212172 3556
rect 212224 3544 212230 3596
rect 251266 3544 251272 3596
rect 251324 3584 251330 3596
rect 252370 3584 252376 3596
rect 251324 3556 252376 3584
rect 251324 3544 251330 3556
rect 252370 3544 252376 3556
rect 252428 3544 252434 3596
rect 259454 3544 259460 3596
rect 259512 3544 259518 3596
rect 103480 3488 104204 3516
rect 103480 3476 103486 3488
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 111886 3516 111892 3528
rect 106976 3488 111892 3516
rect 106976 3476 106982 3488
rect 111886 3476 111892 3488
rect 111944 3476 111950 3528
rect 116118 3476 116124 3528
rect 116176 3516 116182 3528
rect 117590 3516 117596 3528
rect 116176 3488 117596 3516
rect 116176 3476 116182 3488
rect 117590 3476 117596 3488
rect 117648 3476 117654 3528
rect 135898 3476 135904 3528
rect 135956 3516 135962 3528
rect 160094 3516 160100 3528
rect 135956 3488 160100 3516
rect 135956 3476 135962 3488
rect 160094 3476 160100 3488
rect 160152 3476 160158 3528
rect 160848 3516 160876 3544
rect 174262 3516 174268 3528
rect 160848 3488 174268 3516
rect 174262 3476 174268 3488
rect 174320 3476 174326 3528
rect 174538 3476 174544 3528
rect 174596 3516 174602 3528
rect 195606 3516 195612 3528
rect 174596 3488 195612 3516
rect 174596 3476 174602 3488
rect 195606 3476 195612 3488
rect 195664 3476 195670 3528
rect 81802 3448 81808 3460
rect 36044 3352 45324 3380
rect 45526 3420 81808 3448
rect 36044 3340 36050 3352
rect 45526 3312 45554 3420
rect 81802 3408 81808 3420
rect 81860 3408 81866 3460
rect 106826 3448 106832 3460
rect 103440 3420 106832 3448
rect 93946 3340 93952 3392
rect 94004 3380 94010 3392
rect 103440 3380 103468 3420
rect 106826 3408 106832 3420
rect 106884 3408 106890 3460
rect 116026 3408 116032 3460
rect 116084 3448 116090 3460
rect 119890 3448 119896 3460
rect 116084 3420 119896 3448
rect 116084 3408 116090 3420
rect 119890 3408 119896 3420
rect 119948 3408 119954 3460
rect 127158 3408 127164 3460
rect 127216 3448 127222 3460
rect 156598 3448 156604 3460
rect 127216 3420 156604 3448
rect 127216 3408 127222 3420
rect 156598 3408 156604 3420
rect 156656 3408 156662 3460
rect 166350 3408 166356 3460
rect 166408 3448 166414 3460
rect 192018 3448 192024 3460
rect 166408 3420 192024 3448
rect 166408 3408 166414 3420
rect 192018 3408 192024 3420
rect 192076 3408 192082 3460
rect 259472 3448 259500 3544
rect 259564 3516 259592 3624
rect 422938 3612 422944 3664
rect 422996 3652 423002 3664
rect 583386 3652 583392 3664
rect 422996 3624 583392 3652
rect 422996 3612 423002 3624
rect 583386 3612 583392 3624
rect 583444 3612 583450 3664
rect 267734 3544 267740 3596
rect 267792 3584 267798 3596
rect 268470 3584 268476 3596
rect 267792 3556 268476 3584
rect 267792 3544 267798 3556
rect 268470 3544 268476 3556
rect 268528 3544 268534 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 276750 3584 276756 3596
rect 276072 3556 276756 3584
rect 276072 3544 276078 3556
rect 276750 3544 276756 3556
rect 276808 3544 276814 3596
rect 307846 3544 307852 3596
rect 307904 3584 307910 3596
rect 309042 3584 309048 3596
rect 307904 3556 309048 3584
rect 307904 3544 307910 3556
rect 309042 3544 309048 3556
rect 309100 3544 309106 3596
rect 316034 3544 316040 3596
rect 316092 3584 316098 3596
rect 317322 3584 317328 3596
rect 316092 3556 317328 3584
rect 316092 3544 316098 3556
rect 317322 3544 317328 3556
rect 317380 3544 317386 3596
rect 324314 3544 324320 3596
rect 324372 3584 324378 3596
rect 325602 3584 325608 3596
rect 324372 3556 325608 3584
rect 324372 3544 324378 3556
rect 325602 3544 325608 3556
rect 325660 3544 325666 3596
rect 332686 3544 332692 3596
rect 332744 3584 332750 3596
rect 333882 3584 333888 3596
rect 332744 3556 333888 3584
rect 332744 3544 332750 3556
rect 333882 3544 333888 3556
rect 333940 3544 333946 3596
rect 357526 3544 357532 3596
rect 357584 3584 357590 3596
rect 358722 3584 358728 3596
rect 357584 3556 358728 3584
rect 357584 3544 357590 3556
rect 358722 3544 358728 3556
rect 358780 3544 358786 3596
rect 365806 3544 365812 3596
rect 365864 3584 365870 3596
rect 367002 3584 367008 3596
rect 365864 3556 367008 3584
rect 365864 3544 365870 3556
rect 367002 3544 367008 3556
rect 367060 3544 367066 3596
rect 373994 3544 374000 3596
rect 374052 3584 374058 3596
rect 375282 3584 375288 3596
rect 374052 3556 375288 3584
rect 374052 3544 374058 3556
rect 375282 3544 375288 3556
rect 375340 3544 375346 3596
rect 390554 3544 390560 3596
rect 390612 3584 390618 3596
rect 391842 3584 391848 3596
rect 390612 3556 391848 3584
rect 390612 3544 390618 3556
rect 391842 3544 391848 3556
rect 391900 3544 391906 3596
rect 398834 3544 398840 3596
rect 398892 3584 398898 3596
rect 400122 3584 400128 3596
rect 398892 3556 400128 3584
rect 398892 3544 398898 3556
rect 400122 3544 400128 3556
rect 400180 3544 400186 3596
rect 418798 3544 418804 3596
rect 418856 3584 418862 3596
rect 580994 3584 581000 3596
rect 418856 3556 581000 3584
rect 418856 3544 418862 3556
rect 580994 3544 581000 3556
rect 581052 3544 581058 3596
rect 479334 3516 479340 3528
rect 259564 3488 479340 3516
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 481634 3476 481640 3528
rect 481692 3516 481698 3528
rect 482462 3516 482468 3528
rect 481692 3488 482468 3516
rect 481692 3476 481698 3488
rect 482462 3476 482468 3488
rect 482520 3476 482526 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 498194 3476 498200 3528
rect 498252 3516 498258 3528
rect 499022 3516 499028 3528
rect 498252 3488 499028 3516
rect 498252 3476 498258 3488
rect 499022 3476 499028 3488
rect 499080 3476 499086 3528
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 523034 3476 523040 3528
rect 523092 3516 523098 3528
rect 523862 3516 523868 3528
rect 523092 3488 523868 3516
rect 523092 3476 523098 3488
rect 523862 3476 523868 3488
rect 523920 3476 523926 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 556154 3476 556160 3528
rect 556212 3516 556218 3528
rect 556982 3516 556988 3528
rect 556212 3488 556988 3516
rect 556212 3476 556218 3488
rect 556982 3476 556988 3488
rect 557040 3476 557046 3528
rect 572714 3476 572720 3528
rect 572772 3516 572778 3528
rect 573542 3516 573548 3528
rect 572772 3488 573548 3516
rect 572772 3476 572778 3488
rect 573542 3476 573548 3488
rect 573600 3476 573606 3528
rect 582190 3448 582196 3460
rect 259472 3420 582196 3448
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 94004 3352 103468 3380
rect 94004 3340 94010 3352
rect 423674 3340 423680 3392
rect 423732 3380 423738 3392
rect 424962 3380 424968 3392
rect 423732 3352 424968 3380
rect 423732 3340 423738 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 432046 3340 432052 3392
rect 432104 3380 432110 3392
rect 433242 3380 433248 3392
rect 432104 3352 433248 3380
rect 432104 3340 432110 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 26206 3284 45554 3312
rect 96246 3272 96252 3324
rect 96304 3312 96310 3324
rect 103422 3312 103428 3324
rect 96304 3284 103428 3312
rect 96304 3272 96310 3284
rect 103422 3272 103428 3284
rect 103480 3272 103486 3324
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 25498 3040 25504 3052
rect 19484 3012 25504 3040
rect 19484 3000 19490 3012
rect 25498 3000 25504 3012
rect 25556 3000 25562 3052
rect 184198 2932 184204 2984
rect 184256 2972 184262 2984
rect 189718 2972 189724 2984
rect 184256 2944 189724 2972
rect 184256 2932 184262 2944
rect 189718 2932 189724 2944
rect 189776 2932 189782 2984
rect 415394 2864 415400 2916
rect 415452 2904 415458 2916
rect 416682 2904 416688 2916
rect 415452 2876 416688 2904
rect 415452 2864 415458 2876
rect 416682 2864 416688 2876
rect 416740 2864 416746 2916
rect 299474 2728 299480 2780
rect 299532 2768 299538 2780
rect 300762 2768 300768 2780
rect 299532 2740 300768 2768
rect 299532 2728 299538 2740
rect 300762 2728 300768 2740
rect 300820 2728 300826 2780
rect 407114 2592 407120 2644
rect 407172 2632 407178 2644
rect 408402 2632 408408 2644
rect 407172 2604 408408 2632
rect 407172 2592 407178 2604
rect 408402 2592 408408 2604
rect 408460 2592 408466 2644
rect 340874 2320 340880 2372
rect 340932 2360 340938 2372
rect 342162 2360 342168 2372
rect 340932 2332 342168 2360
rect 340932 2320 340938 2332
rect 342162 2320 342168 2332
rect 342220 2320 342226 2372
rect 349154 2320 349160 2372
rect 349212 2360 349218 2372
rect 350442 2360 350448 2372
rect 349212 2332 350448 2360
rect 349212 2320 349218 2332
rect 350442 2320 350448 2332
rect 350500 2320 350506 2372
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 170312 700544 170364 700596
rect 180064 700544 180116 700596
rect 105452 700476 105504 700528
rect 185584 700476 185636 700528
rect 535736 700476 535788 700528
rect 543464 700476 543516 700528
rect 89168 700408 89220 700460
rect 543004 700408 543056 700460
rect 24308 700340 24360 700392
rect 543832 700340 543884 700392
rect 8116 700272 8168 700324
rect 543924 700272 543976 700324
rect 348792 700068 348844 700120
rect 349804 700068 349856 700120
rect 218980 699660 219032 699712
rect 220084 699660 220136 699712
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 534356 696940 534408 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 193864 683136 193916 683188
rect 535552 683136 535604 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 545304 670692 545356 670744
rect 3424 656888 3476 656940
rect 545212 656888 545264 656940
rect 554044 643084 554096 643136
rect 580172 643084 580224 643136
rect 534172 630640 534224 630692
rect 579988 630640 580040 630692
rect 3516 618264 3568 618316
rect 544384 618264 544436 618316
rect 533344 616836 533396 616888
rect 580172 616836 580224 616888
rect 3516 605820 3568 605872
rect 546776 605820 546828 605872
rect 153200 599564 153252 599616
rect 542636 599564 542688 599616
rect 532884 590656 532936 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 202880 579640 202932 579692
rect 546592 579640 546644 579692
rect 532792 576852 532844 576904
rect 580172 576852 580224 576904
rect 3240 565836 3292 565888
rect 177304 565836 177356 565888
rect 3332 553392 3384 553444
rect 546684 553392 546736 553444
rect 2964 527144 3016 527196
rect 208400 527144 208452 527196
rect 548156 527144 548208 527196
rect 531320 524424 531372 524476
rect 580172 524424 580224 524476
rect 3516 514768 3568 514820
rect 177396 514768 177448 514820
rect 299480 511912 299532 511964
rect 300124 511912 300176 511964
rect 300124 510620 300176 510672
rect 539876 510620 539928 510672
rect 3056 500964 3108 501016
rect 547972 500964 548024 501016
rect 477500 497496 477552 497548
rect 536840 497496 536892 497548
rect 282920 497428 282972 497480
rect 539692 497428 539744 497480
rect 530124 484372 530176 484424
rect 580172 484372 580224 484424
rect 531412 470568 531464 470620
rect 579988 470568 580040 470620
rect 530584 456764 530636 456816
rect 580172 456764 580224 456816
rect 527180 453296 527232 453348
rect 535644 453296 535696 453348
rect 529664 430584 529716 430636
rect 580172 430584 580224 430636
rect 412640 428748 412692 428800
rect 538496 428748 538548 428800
rect 349804 428680 349856 428732
rect 539784 428816 539836 428868
rect 220084 428612 220136 428664
rect 541532 428748 541584 428800
rect 539692 428612 539744 428664
rect 540520 428612 540572 428664
rect 177396 428544 177448 428596
rect 548892 428544 548944 428596
rect 177304 428476 177356 428528
rect 548064 428476 548116 428528
rect 3608 428408 3660 428460
rect 549996 428408 550048 428460
rect 534356 427456 534408 427508
rect 554044 427456 554096 427508
rect 531872 427388 531924 427440
rect 580448 427388 580500 427440
rect 462320 427320 462372 427372
rect 537024 427320 537076 427372
rect 397460 427252 397512 427304
rect 538220 427252 538272 427304
rect 201500 427184 201552 427236
rect 541164 427184 541216 427236
rect 71780 427116 71832 427168
rect 543280 427116 543332 427168
rect 3700 427048 3752 427100
rect 549628 427048 549680 427100
rect 364340 426368 364392 426420
rect 364984 426368 365036 426420
rect 535184 425892 535236 425944
rect 580264 425892 580316 425944
rect 331220 425824 331272 425876
rect 539140 425824 539192 425876
rect 3516 425756 3568 425808
rect 212540 425756 212592 425808
rect 266360 425756 266412 425808
rect 540152 425756 540204 425808
rect 136640 425688 136692 425740
rect 542360 425688 542412 425740
rect 184940 425552 184992 425604
rect 185584 425552 185636 425604
rect 364984 425212 365036 425264
rect 538864 425212 538916 425264
rect 212540 425144 212592 425196
rect 549352 425144 549404 425196
rect 185584 425076 185636 425128
rect 543096 425076 543148 425128
rect 234620 425008 234672 425060
rect 235264 425008 235316 425060
rect 543004 425008 543056 425060
rect 543740 425008 543792 425060
rect 532792 424668 532844 424720
rect 533160 424668 533212 424720
rect 445024 424396 445076 424448
rect 494060 424600 494112 424652
rect 536840 424600 536892 424652
rect 536748 424532 536800 424584
rect 558920 424532 558972 424584
rect 532792 424464 532844 424516
rect 580356 424464 580408 424516
rect 531688 424396 531740 424448
rect 580540 424396 580592 424448
rect 3424 424328 3476 424380
rect 198740 424328 198792 424380
rect 429200 424328 429252 424380
rect 529204 424328 529256 424380
rect 235264 423920 235316 423972
rect 540980 423920 541032 423972
rect 198740 423852 198792 423904
rect 544384 423920 544436 423972
rect 546960 423920 547012 423972
rect 546132 423852 546184 423904
rect 546684 423852 546736 423904
rect 547512 423852 547564 423904
rect 179420 423784 179472 423836
rect 180064 423784 180116 423836
rect 541900 423784 541952 423836
rect 543832 423784 543884 423836
rect 544752 423784 544804 423836
rect 546592 423784 546644 423836
rect 547144 423784 547196 423836
rect 547972 423784 548024 423836
rect 548616 423784 548668 423836
rect 77944 423716 77996 423768
rect 556988 423716 557040 423768
rect 4896 423648 4948 423700
rect 530124 423580 530176 423632
rect 530860 423580 530912 423632
rect 531320 423580 531372 423632
rect 532056 423580 532108 423632
rect 550364 423512 550416 423564
rect 445300 423240 445352 423292
rect 533528 423240 533580 423292
rect 445116 423172 445168 423224
rect 535736 423172 535788 423224
rect 536748 423172 536800 423224
rect 524144 423104 524196 423156
rect 547788 423104 547840 423156
rect 175924 423036 175976 423088
rect 553584 423036 553636 423088
rect 4068 422968 4120 423020
rect 4896 422968 4948 423020
rect 87604 422968 87656 423020
rect 552204 422968 552256 423020
rect 43444 422900 43496 422952
rect 551008 422900 551060 422952
rect 522948 422832 523000 422884
rect 549260 422832 549312 422884
rect 522028 422764 522080 422816
rect 561036 422764 561088 422816
rect 529020 422696 529072 422748
rect 548524 422696 548576 422748
rect 445208 422628 445260 422680
rect 534724 422628 534776 422680
rect 535184 422628 535236 422680
rect 535276 422628 535328 422680
rect 558368 422628 558420 422680
rect 530492 422560 530544 422612
rect 561680 422560 561732 422612
rect 352564 422492 352616 422544
rect 554228 422492 554280 422544
rect 525708 422424 525760 422476
rect 535368 422424 535420 422476
rect 526260 422356 526312 422408
rect 538772 422356 538824 422408
rect 523776 422288 523828 422340
rect 529940 422288 529992 422340
rect 550640 422288 550692 422340
rect 558092 422288 558144 422340
rect 126980 421948 127032 422000
rect 530768 421948 530820 422000
rect 284944 421880 284996 421932
rect 529296 421880 529348 421932
rect 548524 421880 548576 421932
rect 580816 421880 580868 421932
rect 527640 421812 527692 421864
rect 560668 421812 560720 421864
rect 528468 421744 528520 421796
rect 560760 421744 560812 421796
rect 136640 421676 136692 421728
rect 532792 421676 532844 421728
rect 535368 421676 535420 421728
rect 580724 421676 580776 421728
rect 3700 421608 3752 421660
rect 527088 421608 527140 421660
rect 529940 421608 529992 421660
rect 580540 421608 580592 421660
rect 3884 421540 3936 421592
rect 550640 421540 550692 421592
rect 528928 421472 528980 421524
rect 563888 421472 563940 421524
rect 528008 421404 528060 421456
rect 563796 421404 563848 421456
rect 526904 421336 526956 421388
rect 562416 421336 562468 421388
rect 521016 421268 521068 421320
rect 560944 421268 560996 421320
rect 521568 421200 521620 421252
rect 561128 421200 561180 421252
rect 520648 421132 520700 421184
rect 580264 421132 580316 421184
rect 522764 421064 522816 421116
rect 561220 421064 561272 421116
rect 524880 420996 524932 421048
rect 562324 420996 562376 421048
rect 525248 420928 525300 420980
rect 569224 420928 569276 420980
rect 529204 420860 529256 420912
rect 537668 420860 537720 420912
rect 538772 420588 538824 420640
rect 542728 420588 542780 420640
rect 525892 420452 525944 420504
rect 539416 420452 539468 420504
rect 524512 420384 524564 420436
rect 541348 420384 541400 420436
rect 541624 420384 541676 420436
rect 547972 420384 548024 420436
rect 549260 420384 549312 420436
rect 580356 420384 580408 420436
rect 530124 420316 530176 420368
rect 546684 420316 546736 420368
rect 547788 420316 547840 420368
rect 580448 420316 580500 420368
rect 530032 420248 530084 420300
rect 541624 420248 541676 420300
rect 542728 420248 542780 420300
rect 580632 420248 580684 420300
rect 232504 420180 232556 420232
rect 553676 420180 553728 420232
rect 132500 420112 132552 420164
rect 531688 420112 531740 420164
rect 539416 420112 539468 420164
rect 546592 420112 546644 420164
rect 160100 420044 160152 420096
rect 429200 420044 429252 420096
rect 529480 420044 529532 420096
rect 562508 420044 562560 420096
rect 527364 419976 527416 420028
rect 445484 419840 445536 419892
rect 530032 419908 530084 419960
rect 541348 419976 541400 420028
rect 560392 419976 560444 420028
rect 445668 419772 445720 419824
rect 525892 419772 525944 419824
rect 236644 419704 236696 419756
rect 530124 419840 530176 419892
rect 528376 419772 528428 419824
rect 193864 419636 193916 419688
rect 519820 419568 519872 419620
rect 193220 419500 193272 419552
rect 193864 419500 193916 419552
rect 514668 419500 514720 419552
rect 517520 419500 517572 419552
rect 545212 419772 545264 419824
rect 519820 418956 519872 419008
rect 547972 419840 548024 419892
rect 555700 419908 555752 419960
rect 546592 419772 546644 419824
rect 546684 419772 546736 419824
rect 554596 419772 554648 419824
rect 556712 419772 556764 419824
rect 559288 419772 559340 419824
rect 559932 419772 559984 419824
rect 560024 419772 560076 419824
rect 560208 419772 560260 419824
rect 563704 419568 563756 419620
rect 566464 419500 566516 419552
rect 561680 419432 561732 419484
rect 580172 419432 580224 419484
rect 447600 416848 447652 416900
rect 517520 416848 517572 416900
rect 447876 416780 447928 416832
rect 517612 416780 517664 416832
rect 448980 415420 449032 415472
rect 517520 415420 517572 415472
rect 449072 413992 449124 414044
rect 517520 413992 517572 414044
rect 450360 412632 450412 412684
rect 517520 412632 517572 412684
rect 450268 411272 450320 411324
rect 517520 411272 517572 411324
rect 3332 411204 3384 411256
rect 43444 411204 43496 411256
rect 447692 409844 447744 409896
rect 517520 409844 517572 409896
rect 450176 408484 450228 408536
rect 517520 408484 517572 408536
rect 449992 407192 450044 407244
rect 517520 407192 517572 407244
rect 450084 407124 450136 407176
rect 517612 407124 517664 407176
rect 449900 405696 449952 405748
rect 517520 405696 517572 405748
rect 562508 405628 562560 405680
rect 580172 405628 580224 405680
rect 447784 404336 447836 404388
rect 517520 404336 517572 404388
rect 449164 402976 449216 403028
rect 517704 402976 517756 403028
rect 449348 401616 449400 401668
rect 517704 401616 517756 401668
rect 449532 400256 449584 400308
rect 517704 400256 517756 400308
rect 449256 400188 449308 400240
rect 517796 400188 517848 400240
rect 449624 398828 449676 398880
rect 517704 398828 517756 398880
rect 449440 397468 449492 397520
rect 517704 397468 517756 397520
rect 449716 396040 449768 396092
rect 517704 396040 517756 396092
rect 450820 394748 450872 394800
rect 517704 394748 517756 394800
rect 449808 394680 449860 394732
rect 517796 394680 517848 394732
rect 447048 393320 447100 393372
rect 517704 393320 517756 393372
rect 448152 392096 448204 392148
rect 517704 392096 517756 392148
rect 447968 392028 448020 392080
rect 517888 392028 517940 392080
rect 446956 391960 447008 392012
rect 517980 391960 518032 392012
rect 448060 390600 448112 390652
rect 517704 390600 517756 390652
rect 446864 390532 446916 390584
rect 517888 390532 517940 390584
rect 448244 389240 448296 389292
rect 517704 389240 517756 389292
rect 446772 389172 446824 389224
rect 517888 389172 517940 389224
rect 448336 387948 448388 388000
rect 517888 387948 517940 388000
rect 446680 387880 446732 387932
rect 517704 387880 517756 387932
rect 446588 387812 446640 387864
rect 517980 387812 518032 387864
rect 448428 386452 448480 386504
rect 517888 386452 517940 386504
rect 446496 386384 446548 386436
rect 517704 386384 517756 386436
rect 517612 379856 517664 379908
rect 550640 379856 550692 379908
rect 563888 379448 563940 379500
rect 580172 379448 580224 379500
rect 519360 379108 519412 379160
rect 549628 379108 549680 379160
rect 519084 379040 519136 379092
rect 549720 379040 549772 379092
rect 518992 378972 519044 379024
rect 549812 378972 549864 379024
rect 519452 378904 519504 378956
rect 550732 378904 550784 378956
rect 519176 378836 519228 378888
rect 550824 378836 550876 378888
rect 519268 378768 519320 378820
rect 550916 378768 550968 378820
rect 521568 378020 521620 378072
rect 523040 378020 523092 378072
rect 521292 377680 521344 377732
rect 533344 377680 533396 377732
rect 524328 377612 524380 377664
rect 549904 377612 549956 377664
rect 523408 377544 523460 377596
rect 549996 377544 550048 377596
rect 524052 377476 524104 377528
rect 551468 377476 551520 377528
rect 520372 377408 520424 377460
rect 549260 377408 549312 377460
rect 524696 376116 524748 376168
rect 550088 376116 550140 376168
rect 523132 376048 523184 376100
rect 551284 376048 551336 376100
rect 523040 375980 523092 376032
rect 552112 375980 552164 376032
rect 523776 374756 523828 374808
rect 551376 374756 551428 374808
rect 520648 374688 520700 374740
rect 551192 374688 551244 374740
rect 520096 374620 520148 374672
rect 551100 374620 551152 374672
rect 533344 371900 533396 371952
rect 552020 371900 552072 371952
rect 521016 371832 521068 371884
rect 549352 371832 549404 371884
rect 3332 371220 3384 371272
rect 222200 371220 222252 371272
rect 223488 371220 223540 371272
rect 522856 371152 522908 371204
rect 552480 371152 552532 371204
rect 522488 371084 522540 371136
rect 552388 371084 552440 371136
rect 522212 371016 522264 371068
rect 552296 371016 552348 371068
rect 521936 370948 521988 371000
rect 552204 370948 552256 371000
rect 518900 370880 518952 370932
rect 549536 370880 549588 370932
rect 517520 370812 517572 370864
rect 549444 370812 549496 370864
rect 518256 370744 518308 370796
rect 551008 370744 551060 370796
rect 518716 370676 518768 370728
rect 553584 370676 553636 370728
rect 518808 370608 518860 370660
rect 553676 370608 553728 370660
rect 514668 370540 514720 370592
rect 553768 370540 553820 370592
rect 450728 370472 450780 370524
rect 518164 370472 518216 370524
rect 518624 370472 518676 370524
rect 553492 370472 553544 370524
rect 3056 358708 3108 358760
rect 87604 358708 87656 358760
rect 560760 353200 560812 353252
rect 579620 353200 579672 353252
rect 549904 352520 549956 352572
rect 560760 352520 560812 352572
rect 2964 346332 3016 346384
rect 444748 346332 444800 346384
rect 563796 325592 563848 325644
rect 580172 325592 580224 325644
rect 226340 320084 226392 320136
rect 226984 320084 227036 320136
rect 3332 319404 3384 319456
rect 226340 319404 226392 319456
rect 566464 313216 566516 313268
rect 580172 313216 580224 313268
rect 3332 306280 3384 306332
rect 175924 306280 175976 306332
rect 561588 299412 561640 299464
rect 580172 299412 580224 299464
rect 113180 298732 113232 298784
rect 560668 298732 560720 298784
rect 561588 298732 561640 298784
rect 446496 298052 446548 298104
rect 460756 298052 460808 298104
rect 545212 298052 545264 298104
rect 553400 298052 553452 298104
rect 450820 297984 450872 298036
rect 482652 297984 482704 298036
rect 535828 297984 535880 298036
rect 553492 297984 553544 298036
rect 446956 297916 447008 297968
rect 476396 297916 476448 297968
rect 538956 297916 539008 297968
rect 553584 297916 553636 297968
rect 446864 297848 446916 297900
rect 473268 297848 473320 297900
rect 542084 297848 542136 297900
rect 553676 297848 553728 297900
rect 446772 297780 446824 297832
rect 470140 297780 470192 297832
rect 510804 297780 510856 297832
rect 550916 297780 550968 297832
rect 446588 297712 446640 297764
rect 467012 297712 467064 297764
rect 513932 297712 513984 297764
rect 549812 297712 549864 297764
rect 446680 297644 446732 297696
rect 463884 297644 463936 297696
rect 517060 297644 517112 297696
rect 550640 297644 550692 297696
rect 447048 297576 447100 297628
rect 479524 297576 479576 297628
rect 520188 297576 520240 297628
rect 549536 297576 549588 297628
rect 523316 297508 523368 297560
rect 551008 297508 551060 297560
rect 498292 297440 498344 297492
rect 550732 297440 550784 297492
rect 501420 297372 501472 297424
rect 549628 297372 549680 297424
rect 504548 297304 504600 297356
rect 550824 297304 550876 297356
rect 507676 297236 507728 297288
rect 549720 297236 549772 297288
rect 526444 297168 526496 297220
rect 549444 297168 549496 297220
rect 3240 293904 3292 293956
rect 444932 293904 444984 293956
rect 562416 273164 562468 273216
rect 580172 273164 580224 273216
rect 231860 267180 231912 267232
rect 232504 267180 232556 267232
rect 3332 266976 3384 267028
rect 231860 266976 231912 267028
rect 563704 259360 563756 259412
rect 579804 259360 579856 259412
rect 2964 255212 3016 255264
rect 352564 255212 352616 255264
rect 560576 245556 560628 245608
rect 580172 245556 580224 245608
rect 440884 244876 440936 244928
rect 560576 244876 560628 244928
rect 109040 224204 109092 224256
rect 440884 224204 440936 224256
rect 3332 214548 3384 214600
rect 236000 214548 236052 214600
rect 236644 214548 236696 214600
rect 560484 206932 560536 206984
rect 579804 206932 579856 206984
rect 103980 206252 104032 206304
rect 560484 206252 560536 206304
rect 170312 203736 170364 203788
rect 300124 203736 300176 203788
rect 40040 203668 40092 203720
rect 189080 203668 189132 203720
rect 165620 203600 165672 203652
rect 364984 203600 365036 203652
rect 4896 203532 4948 203584
rect 218152 203532 218204 203584
rect 189080 202784 189132 202836
rect 189724 202784 189776 202836
rect 445392 202784 445444 202836
rect 123668 202512 123720 202564
rect 284944 202512 284996 202564
rect 156880 202444 156932 202496
rect 445024 202444 445076 202496
rect 152096 202376 152148 202428
rect 445116 202376 445168 202428
rect 147404 202308 147456 202360
rect 445208 202308 445260 202360
rect 142620 202240 142672 202292
rect 445300 202240 445352 202292
rect 175832 202172 175884 202224
rect 235264 202172 235316 202224
rect 256056 202172 256108 202224
rect 559932 202172 559984 202224
rect 118976 202104 119028 202156
rect 549904 202104 549956 202156
rect 100024 201628 100076 201680
rect 261576 201628 261628 201680
rect 95148 201560 95200 201612
rect 260104 201560 260156 201612
rect 3792 201492 3844 201544
rect 256056 201492 256108 201544
rect 561312 201424 561364 201476
rect 564440 201424 564492 201476
rect 251364 200880 251416 200932
rect 445576 200880 445628 200932
rect 246580 200812 246632 200864
rect 445668 200812 445720 200864
rect 241888 200744 241940 200796
rect 445484 200744 445536 200796
rect 85488 200472 85540 200524
rect 261484 200472 261536 200524
rect 4896 200404 4948 200456
rect 241888 200404 241940 200456
rect 3884 200336 3936 200388
rect 246580 200336 246632 200388
rect 3700 200268 3752 200320
rect 251364 200268 251416 200320
rect 90548 200200 90600 200252
rect 438124 200200 438176 200252
rect 81072 200132 81124 200184
rect 561312 200132 561364 200184
rect 562324 193128 562376 193180
rect 579620 193128 579672 193180
rect 569224 179324 569276 179376
rect 579620 179324 579672 179376
rect 261576 166948 261628 167000
rect 560392 166948 560444 167000
rect 580172 166948 580224 167000
rect 2780 162936 2832 162988
rect 4896 162936 4948 162988
rect 2780 150152 2832 150204
rect 4988 150152 5040 150204
rect 3516 137912 3568 137964
rect 79324 137912 79376 137964
rect 260104 126896 260156 126948
rect 560024 126896 560076 126948
rect 580172 126896 580224 126948
rect 561220 113092 561272 113144
rect 579620 113092 579672 113144
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 438124 86912 438176 86964
rect 560300 86844 560352 86896
rect 580172 86912 580224 86964
rect 2964 85484 3016 85536
rect 77944 85484 77996 85536
rect 80750 79840 80802 79892
rect 89812 79840 89864 79892
rect 90686 79840 90738 79892
rect 96712 79840 96764 79892
rect 97586 79840 97638 79892
rect 98092 79840 98144 79892
rect 99058 79840 99110 79892
rect 121552 79840 121604 79892
rect 122426 79840 122478 79892
rect 123530 79840 123582 79892
rect 80060 79772 80112 79824
rect 80152 79772 80204 79824
rect 81118 79772 81170 79824
rect 81624 79772 81676 79824
rect 82222 79772 82274 79824
rect 89720 79772 89772 79824
rect 90318 79772 90370 79824
rect 96620 79772 96672 79824
rect 97218 79772 97270 79824
rect 98184 79772 98236 79824
rect 98690 79772 98742 79824
rect 99564 79772 99616 79824
rect 100530 79772 100582 79824
rect 103612 79772 103664 79824
rect 104486 79772 104538 79824
rect 106372 79772 106424 79824
rect 107062 79772 107114 79824
rect 111984 79772 112036 79824
rect 112582 79772 112634 79824
rect 116032 79772 116084 79824
rect 116906 79772 116958 79824
rect 121460 79772 121512 79824
rect 122058 79772 122110 79824
rect 79968 79636 80020 79688
rect 80244 79636 80296 79688
rect 122840 79636 122892 79688
rect 139998 79840 140050 79892
rect 146300 79840 146352 79892
rect 147266 79840 147318 79892
rect 151820 79840 151872 79892
rect 152694 79840 152746 79892
rect 157340 79840 157392 79892
rect 157846 79840 157898 79892
rect 158214 79840 158266 79892
rect 124312 79772 124364 79824
rect 125370 79772 125422 79824
rect 126980 79772 127032 79824
rect 128222 79772 128274 79824
rect 129924 79772 129976 79824
rect 130798 79772 130850 79824
rect 132500 79772 132552 79824
rect 133006 79772 133058 79824
rect 133972 79772 134024 79824
rect 134846 79772 134898 79824
rect 139584 79772 139636 79824
rect 140780 79772 140832 79824
rect 141746 79772 141798 79824
rect 144920 79772 144972 79824
rect 146162 79772 146214 79824
rect 146392 79772 146444 79824
rect 146898 79772 146950 79824
rect 147864 79772 147916 79824
rect 148738 79772 148790 79824
rect 152004 79772 152056 79824
rect 153062 79772 153114 79824
rect 153200 79772 153252 79824
rect 154166 79772 154218 79824
rect 156144 79772 156196 79824
rect 157110 79772 157162 79824
rect 157432 79636 157484 79688
rect 170634 79840 170686 79892
rect 162860 79772 162912 79824
rect 163734 79772 163786 79824
rect 164240 79772 164292 79824
rect 164746 79772 164798 79824
rect 167000 79772 167052 79824
rect 168058 79772 168110 79824
rect 169852 79772 169904 79824
rect 171232 79772 171284 79824
rect 172106 79772 172158 79824
rect 174314 79840 174366 79892
rect 174682 79840 174734 79892
rect 183652 79840 183704 79892
rect 184526 79840 184578 79892
rect 189080 79840 189132 79892
rect 189954 79840 190006 79892
rect 200534 79840 200586 79892
rect 200902 79840 200954 79892
rect 206422 79840 206474 79892
rect 173900 79636 173952 79688
rect 173992 79636 174044 79688
rect 176660 79772 176712 79824
rect 177534 79772 177586 79824
rect 178040 79772 178092 79824
rect 178638 79772 178690 79824
rect 182180 79772 182232 79824
rect 183054 79772 183106 79824
rect 183560 79772 183612 79824
rect 184158 79772 184210 79824
rect 187792 79772 187844 79824
rect 188850 79772 188902 79824
rect 190460 79772 190512 79824
rect 191058 79772 191110 79824
rect 193404 79772 193456 79824
rect 194370 79772 194422 79824
rect 194600 79772 194652 79824
rect 195474 79772 195526 79824
rect 198924 79772 198976 79824
rect 199890 79772 199942 79824
rect 200120 79636 200172 79688
rect 200212 79636 200264 79688
rect 204352 79772 204404 79824
rect 205318 79772 205370 79824
rect 205640 79636 205692 79688
rect 225374 79840 225426 79892
rect 229790 79840 229842 79892
rect 230894 79840 230946 79892
rect 231262 79840 231314 79892
rect 231860 79840 231912 79892
rect 232366 79840 232418 79892
rect 232734 79840 232786 79892
rect 208400 79772 208452 79824
rect 208998 79772 209050 79824
rect 209780 79772 209832 79824
rect 210838 79772 210890 79824
rect 213920 79772 213972 79824
rect 215162 79772 215214 79824
rect 219440 79772 219492 79824
rect 219946 79772 219998 79824
rect 220912 79772 220964 79824
rect 221786 79772 221838 79824
rect 222292 79772 222344 79824
rect 223258 79772 223310 79824
rect 224960 79772 225012 79824
rect 225052 79772 225104 79824
rect 226110 79772 226162 79824
rect 227720 79772 227772 79824
rect 228686 79772 228738 79824
rect 229100 79772 229152 79824
rect 224868 79636 224920 79688
rect 225236 79636 225288 79688
rect 230480 79636 230532 79688
rect 230572 79636 230624 79688
rect 231952 79636 232004 79688
rect 238162 79840 238214 79892
rect 244280 79840 244332 79892
rect 244786 79840 244838 79892
rect 248748 79840 248800 79892
rect 249616 79840 249668 79892
rect 251180 79840 251232 79892
rect 251686 79840 251738 79892
rect 252652 79840 252704 79892
rect 253526 79840 253578 79892
rect 254124 79840 254176 79892
rect 254998 79840 255050 79892
rect 238760 79772 238812 79824
rect 239634 79772 239686 79824
rect 241704 79772 241756 79824
rect 242578 79772 242630 79824
rect 248420 79772 248472 79824
rect 249110 79772 249162 79824
rect 252560 79772 252612 79824
rect 253158 79772 253210 79824
rect 254032 79772 254084 79824
rect 254630 79772 254682 79824
rect 256792 79772 256844 79824
rect 257942 79772 257994 79824
rect 258080 79772 258132 79824
rect 258678 79772 258730 79824
rect 237380 79636 237432 79688
rect 80336 78752 80388 78804
rect 447784 78752 447836 78804
rect 80244 78684 80296 78736
rect 447876 78684 447928 78736
rect 112168 78616 112220 78668
rect 114560 78616 114612 78668
rect 189632 78616 189684 78668
rect 191380 78616 191432 78668
rect 97264 78548 97316 78600
rect 105268 78548 105320 78600
rect 188528 78548 188580 78600
rect 192576 78548 192628 78600
rect 70400 78480 70452 78532
rect 101956 78480 102008 78532
rect 131580 78480 131632 78532
rect 134524 78480 134576 78532
rect 185676 78480 185728 78532
rect 191288 78480 191340 78532
rect 204996 78480 205048 78532
rect 210424 78480 210476 78532
rect 65524 78412 65576 78464
rect 99748 78412 99800 78464
rect 53104 78344 53156 78396
rect 93216 78344 93268 78396
rect 110420 78344 110472 78396
rect 114008 78344 114060 78396
rect 50344 78276 50396 78328
rect 91100 78276 91152 78328
rect 93124 78276 93176 78328
rect 96436 78276 96488 78328
rect 227996 78276 228048 78328
rect 258724 78276 258776 78328
rect 28264 78208 28316 78260
rect 86224 78208 86276 78260
rect 110512 78208 110564 78260
rect 111064 78208 111116 78260
rect 207204 78208 207256 78260
rect 213092 78208 213144 78260
rect 226892 78208 226944 78260
rect 289084 78208 289136 78260
rect 32404 78140 32456 78192
rect 88800 78140 88852 78192
rect 136364 78140 136416 78192
rect 166448 78140 166500 78192
rect 215944 78140 215996 78192
rect 226984 78140 227036 78192
rect 259092 78140 259144 78192
rect 418804 78140 418856 78192
rect 25504 78072 25556 78124
rect 85948 78072 86000 78124
rect 101404 78072 101456 78124
rect 106280 78072 106332 78124
rect 111064 78072 111116 78124
rect 113640 78072 113692 78124
rect 129372 78072 129424 78124
rect 135904 78072 135956 78124
rect 153844 78072 153896 78124
rect 188344 78072 188396 78124
rect 209412 78072 209464 78124
rect 214564 78072 214616 78124
rect 220360 78072 220412 78124
rect 255964 78072 256016 78124
rect 260104 78072 260156 78124
rect 422944 78072 422996 78124
rect 15844 78004 15896 78056
rect 83280 78004 83332 78056
rect 120632 78004 120684 78056
rect 126244 78004 126296 78056
rect 149520 78004 149572 78056
rect 187056 78004 187108 78056
rect 198464 78004 198516 78056
rect 203524 78004 203576 78056
rect 208308 78004 208360 78056
rect 213184 78004 213236 78056
rect 222568 78004 222620 78056
rect 407764 78004 407816 78056
rect 10324 77936 10376 77988
rect 81440 77936 81492 77988
rect 102140 77936 102192 77988
rect 111800 77936 111852 77988
rect 131948 77936 132000 77988
rect 141424 77936 141476 77988
rect 144000 77936 144052 77988
rect 186964 77936 187016 77988
rect 224684 77936 224736 77988
rect 411904 77936 411956 77988
rect 124220 77868 124272 77920
rect 129096 77868 129148 77920
rect 107660 77800 107712 77852
rect 113272 77800 113324 77852
rect 121368 77800 121420 77852
rect 123484 77800 123536 77852
rect 118424 77732 118476 77784
rect 124220 77732 124272 77784
rect 190736 77664 190788 77716
rect 192392 77664 192444 77716
rect 106924 77460 106976 77512
rect 108856 77460 108908 77512
rect 105544 77392 105596 77444
rect 107384 77392 107436 77444
rect 135628 77392 135680 77444
rect 144184 77460 144236 77512
rect 201684 77460 201736 77512
rect 209044 77460 209096 77512
rect 142436 77392 142488 77444
rect 187516 77392 187568 77444
rect 191104 77392 191156 77444
rect 202788 77392 202840 77444
rect 207756 77392 207808 77444
rect 229192 77392 229244 77444
rect 100024 77324 100076 77376
rect 103060 77324 103112 77376
rect 107016 77324 107068 77376
rect 108488 77324 108540 77376
rect 118056 77324 118108 77376
rect 119344 77324 119396 77376
rect 123208 77324 123260 77376
rect 129004 77324 129056 77376
rect 135352 77324 135404 77376
rect 137284 77324 137336 77376
rect 81532 77256 81584 77308
rect 82544 77256 82596 77308
rect 82912 77256 82964 77308
rect 84016 77256 84068 77308
rect 86960 77256 87012 77308
rect 87236 77256 87288 77308
rect 88524 77256 88576 77308
rect 89536 77256 89588 77308
rect 93952 77256 94004 77308
rect 94136 77256 94188 77308
rect 100852 77256 100904 77308
rect 101588 77256 101640 77308
rect 104992 77256 105044 77308
rect 105912 77256 105964 77308
rect 107752 77256 107804 77308
rect 108120 77256 108172 77308
rect 108304 77256 108356 77308
rect 109592 77256 109644 77308
rect 109684 77256 109736 77308
rect 110696 77256 110748 77308
rect 111892 77256 111944 77308
rect 112904 77256 112956 77308
rect 118792 77256 118844 77308
rect 119804 77256 119856 77308
rect 121000 77256 121052 77308
rect 122104 77256 122156 77308
rect 125784 77256 125836 77308
rect 126428 77256 126480 77308
rect 127992 77256 128044 77308
rect 129188 77256 129240 77308
rect 129740 77256 129792 77308
rect 130384 77256 130436 77308
rect 132684 77256 132736 77308
rect 133328 77256 133380 77308
rect 136732 77256 136784 77308
rect 137376 77256 137428 77308
rect 138204 77256 138256 77308
rect 139216 77256 139268 77308
rect 139492 77256 139544 77308
rect 140596 77256 140648 77308
rect 93860 77188 93912 77240
rect 94964 77188 95016 77240
rect 109224 77188 109276 77240
rect 109960 77188 110012 77240
rect 125692 77188 125744 77240
rect 126796 77188 126848 77240
rect 132592 77188 132644 77240
rect 133696 77188 133748 77240
rect 136640 77188 136692 77240
rect 137744 77188 137796 77240
rect 138112 77188 138164 77240
rect 138848 77188 138900 77240
rect 87144 77120 87196 77172
rect 87696 77120 87748 77172
rect 92572 77120 92624 77172
rect 93492 77120 93544 77172
rect 93952 77120 94004 77172
rect 94596 77120 94648 77172
rect 110696 77120 110748 77172
rect 111432 77120 111484 77172
rect 167184 77324 167236 77376
rect 169024 77324 169076 77376
rect 192944 77324 192996 77376
rect 193864 77324 193916 77376
rect 194048 77324 194100 77376
rect 195244 77324 195296 77376
rect 206100 77324 206152 77376
rect 209136 77324 209188 77376
rect 210516 77324 210568 77376
rect 217324 77324 217376 77376
rect 143632 77256 143684 77308
rect 144644 77256 144696 77308
rect 145104 77256 145156 77308
rect 145748 77256 145800 77308
rect 147680 77256 147732 77308
rect 148324 77256 148376 77308
rect 149060 77256 149112 77308
rect 150164 77256 150216 77308
rect 150624 77256 150676 77308
rect 151636 77256 151688 77308
rect 154580 77256 154632 77308
rect 155592 77256 155644 77308
rect 155960 77256 156012 77308
rect 156696 77256 156748 77308
rect 168472 77256 168524 77308
rect 169484 77256 169536 77308
rect 175372 77256 175424 77308
rect 176384 77256 176436 77308
rect 191840 77256 191892 77308
rect 192024 77256 192076 77308
rect 193220 77256 193272 77308
rect 193588 77256 193640 77308
rect 194692 77256 194744 77308
rect 195060 77256 195112 77308
rect 198740 77256 198792 77308
rect 199476 77256 199528 77308
rect 203892 77256 203944 77308
rect 206284 77256 206336 77308
rect 211252 77256 211304 77308
rect 211528 77256 211580 77308
rect 212632 77256 212684 77308
rect 213276 77256 213328 77308
rect 213736 77256 213788 77308
rect 215944 77256 215996 77308
rect 218152 77256 218204 77308
rect 218336 77256 218388 77308
rect 219532 77256 219584 77308
rect 220636 77256 220688 77308
rect 223672 77256 223724 77308
rect 223856 77256 223908 77308
rect 226432 77256 226484 77308
rect 227536 77256 227588 77308
rect 150532 77188 150584 77240
rect 151268 77188 151320 77240
rect 168380 77188 168432 77240
rect 169116 77188 169168 77240
rect 211160 77188 211212 77240
rect 211712 77188 211764 77240
rect 214104 77188 214156 77240
rect 214748 77188 214800 77240
rect 218060 77188 218112 77240
rect 219164 77188 219216 77240
rect 223580 77188 223632 77240
rect 224224 77188 224276 77240
rect 226524 77188 226576 77240
rect 227168 77188 227220 77240
rect 242992 77324 243044 77376
rect 244004 77324 244056 77376
rect 234620 77256 234672 77308
rect 235632 77256 235684 77308
rect 236092 77256 236144 77308
rect 236644 77256 236696 77308
rect 238944 77256 238996 77308
rect 239956 77256 240008 77308
rect 240232 77256 240284 77308
rect 241060 77256 241112 77308
rect 241520 77256 241572 77308
rect 242164 77256 242216 77308
rect 243084 77256 243136 77308
rect 243636 77256 243688 77308
rect 244464 77256 244516 77308
rect 245476 77256 245528 77308
rect 245752 77256 245804 77308
rect 246580 77256 246632 77308
rect 247132 77256 247184 77308
rect 247684 77256 247736 77308
rect 248512 77256 248564 77308
rect 249432 77256 249484 77308
rect 249800 77256 249852 77308
rect 250352 77256 250404 77308
rect 251364 77256 251416 77308
rect 252376 77256 252428 77308
rect 229284 77188 229336 77240
rect 236000 77188 236052 77240
rect 237012 77188 237064 77240
rect 242900 77188 242952 77240
rect 243268 77188 243320 77240
rect 247040 77188 247092 77240
rect 248052 77188 248104 77240
rect 191840 77120 191892 77172
rect 192484 77120 192536 77172
rect 218152 77120 218204 77172
rect 218796 77120 218848 77172
rect 142436 77052 142488 77104
rect 255596 77052 255648 77104
rect 256424 77052 256476 77104
rect 170036 76780 170088 76832
rect 291200 76780 291252 76832
rect 216772 76712 216824 76764
rect 441620 76712 441672 76764
rect 217784 76644 217836 76696
rect 445760 76644 445812 76696
rect 51080 76576 51132 76628
rect 95700 76576 95752 76628
rect 225236 76576 225288 76628
rect 469220 76576 469272 76628
rect 49700 76508 49752 76560
rect 95332 76508 95384 76560
rect 257620 76508 257672 76560
rect 574100 76508 574152 76560
rect 86960 75624 87012 75676
rect 88064 75624 88116 75676
rect 168840 75420 168892 75472
rect 287060 75420 287112 75472
rect 195888 75352 195940 75404
rect 374000 75352 374052 75404
rect 214472 75284 214524 75336
rect 434720 75284 434772 75336
rect 215576 75216 215628 75268
rect 438860 75216 438912 75268
rect 37280 75148 37332 75200
rect 91744 75148 91796 75200
rect 161572 75148 161624 75200
rect 162584 75148 162636 75200
rect 162952 75148 163004 75200
rect 164056 75148 164108 75200
rect 164332 75148 164384 75200
rect 165068 75148 165120 75200
rect 176844 75148 176896 75200
rect 177856 75148 177908 75200
rect 180800 75148 180852 75200
rect 181904 75148 181956 75200
rect 182364 75148 182416 75200
rect 183376 75148 183428 75200
rect 249616 75148 249668 75200
rect 546500 75148 546552 75200
rect 160008 75080 160060 75132
rect 160284 75080 160336 75132
rect 179328 75080 179380 75132
rect 179604 75080 179656 75132
rect 184848 75080 184900 75132
rect 185124 75080 185176 75132
rect 160192 75012 160244 75064
rect 160744 75012 160796 75064
rect 179512 75012 179564 75064
rect 180064 75012 180116 75064
rect 185032 75012 185084 75064
rect 185952 75012 186004 75064
rect 167460 74060 167512 74112
rect 284300 74060 284352 74112
rect 212632 73992 212684 74044
rect 431960 73992 432012 74044
rect 239036 73924 239088 73976
rect 514760 73924 514812 73976
rect 243176 73856 243228 73908
rect 527180 73856 527232 73908
rect 247316 73788 247368 73840
rect 540980 73788 541032 73840
rect 561128 73108 561180 73160
rect 579988 73108 580040 73160
rect 166632 72700 166684 72752
rect 280160 72700 280212 72752
rect 196716 72632 196768 72684
rect 378140 72632 378192 72684
rect 211804 72564 211856 72616
rect 427820 72564 427872 72616
rect 243084 72496 243136 72548
rect 529940 72496 529992 72548
rect 247224 72428 247276 72480
rect 539600 72428 539652 72480
rect 165528 71272 165580 71324
rect 276020 71272 276072 71324
rect 207112 71204 207164 71256
rect 414020 71204 414072 71256
rect 209964 71136 210016 71188
rect 420920 71136 420972 71188
rect 211344 71068 211396 71120
rect 423680 71068 423732 71120
rect 255596 71000 255648 71052
rect 571340 71000 571392 71052
rect 164424 69912 164476 69964
rect 273260 69912 273312 69964
rect 197820 69844 197872 69896
rect 382280 69844 382332 69896
rect 203432 69776 203484 69828
rect 398840 69776 398892 69828
rect 204444 69708 204496 69760
rect 402980 69708 403032 69760
rect 254216 69640 254268 69692
rect 564532 69640 564584 69692
rect 163136 68552 163188 68604
rect 269120 68552 269172 68604
rect 199016 68484 199068 68536
rect 385040 68484 385092 68536
rect 200396 68416 200448 68468
rect 391940 68416 391992 68468
rect 202144 68348 202196 68400
rect 396080 68348 396132 68400
rect 251456 68280 251508 68332
rect 556160 68280 556212 68332
rect 162032 67124 162084 67176
rect 266360 67124 266412 67176
rect 189724 67056 189776 67108
rect 357440 67056 357492 67108
rect 194784 66988 194836 67040
rect 371240 66988 371292 67040
rect 200304 66920 200356 66972
rect 389180 66920 389232 66972
rect 250444 66852 250496 66904
rect 553400 66852 553452 66904
rect 160928 65764 160980 65816
rect 262220 65764 262272 65816
rect 186872 65696 186924 65748
rect 346400 65696 346452 65748
rect 187884 65628 187936 65680
rect 349160 65628 349212 65680
rect 92756 65560 92808 65612
rect 189172 65560 189224 65612
rect 353300 65560 353352 65612
rect 247132 65492 247184 65544
rect 542360 65492 542412 65544
rect 92756 65356 92808 65408
rect 160284 64404 160336 64456
rect 259552 64404 259604 64456
rect 183744 64336 183796 64388
rect 335360 64336 335412 64388
rect 185124 64268 185176 64320
rect 339500 64268 339552 64320
rect 185032 64200 185084 64252
rect 342260 64200 342312 64252
rect 238944 64132 238996 64184
rect 517520 64132 517572 64184
rect 169944 63044 169996 63096
rect 293960 63044 294012 63096
rect 179696 62976 179748 63028
rect 324320 62976 324372 63028
rect 181076 62908 181128 62960
rect 328460 62908 328512 62960
rect 182456 62840 182508 62892
rect 332600 62840 332652 62892
rect 117320 62772 117372 62824
rect 117504 62772 117556 62824
rect 238852 62772 238904 62824
rect 514852 62772 514904 62824
rect 176936 61616 176988 61668
rect 314660 61616 314712 61668
rect 178132 61548 178184 61600
rect 317420 61548 317472 61600
rect 179604 61480 179656 61532
rect 321560 61480 321612 61532
rect 194692 61412 194744 61464
rect 372620 61412 372672 61464
rect 229376 61344 229428 61396
rect 485780 61344 485832 61396
rect 561036 60664 561088 60716
rect 580172 60664 580224 60716
rect 174084 60256 174136 60308
rect 303620 60256 303672 60308
rect 174176 60188 174228 60240
rect 307760 60188 307812 60240
rect 175556 60120 175608 60172
rect 310520 60120 310572 60172
rect 247040 60052 247092 60104
rect 543740 60052 543792 60104
rect 149152 59984 149204 60036
rect 223672 59984 223724 60036
rect 258172 59984 258224 60036
rect 576860 59984 576912 60036
rect 169852 58964 169904 59016
rect 292580 58964 292632 59016
rect 171324 58896 171376 58948
rect 296720 58896 296772 58948
rect 225144 58828 225196 58880
rect 471980 58828 472032 58880
rect 253940 58760 253992 58812
rect 563060 58760 563112 58812
rect 254124 58692 254176 58744
rect 565820 58692 565872 58744
rect 255504 58624 255556 58676
rect 569960 58624 570012 58676
rect 92664 58556 92716 58608
rect 92848 58556 92900 58608
rect 168564 57536 168616 57588
rect 285680 57536 285732 57588
rect 168472 57468 168524 57520
rect 289820 57468 289872 57520
rect 223856 57400 223908 57452
rect 465080 57400 465132 57452
rect 244556 57332 244608 57384
rect 534080 57332 534132 57384
rect 245844 57264 245896 57316
rect 538220 57264 538272 57316
rect 248604 57196 248656 57248
rect 545120 57196 545172 57248
rect 165712 56176 165764 56228
rect 278780 56176 278832 56228
rect 167092 56108 167144 56160
rect 282920 56108 282972 56160
rect 221004 56040 221056 56092
rect 456800 56040 456852 56092
rect 240324 55972 240376 56024
rect 520280 55972 520332 56024
rect 241796 55904 241848 55956
rect 523040 55904 523092 55956
rect 242992 55836 243044 55888
rect 531320 55836 531372 55888
rect 164332 54816 164384 54868
rect 276112 54816 276164 54868
rect 218336 54748 218388 54800
rect 447140 54748 447192 54800
rect 237472 54680 237524 54732
rect 509240 54680 509292 54732
rect 237656 54612 237708 54664
rect 513380 54612 513432 54664
rect 238760 54544 238812 54596
rect 516140 54544 516192 54596
rect 256884 54476 256936 54528
rect 572720 54476 572772 54528
rect 163044 53388 163096 53440
rect 267740 53388 267792 53440
rect 162952 53320 163004 53372
rect 271880 53320 271932 53372
rect 214104 53252 214156 53304
rect 436100 53252 436152 53304
rect 233424 53184 233476 53236
rect 498200 53184 498252 53236
rect 234896 53116 234948 53168
rect 502340 53116 502392 53168
rect 236276 53048 236328 53100
rect 506480 53048 506532 53100
rect 153292 52028 153344 52080
rect 237472 52028 237524 52080
rect 161664 51960 161716 52012
rect 264980 51960 265032 52012
rect 171232 51892 171284 51944
rect 298100 51892 298152 51944
rect 226524 51824 226576 51876
rect 476120 51824 476172 51876
rect 232044 51756 232096 51808
rect 491300 51756 491352 51808
rect 232136 51688 232188 51740
rect 495440 51688 495492 51740
rect 152096 50668 152148 50720
rect 234896 50668 234948 50720
rect 160192 50600 160244 50652
rect 260840 50600 260892 50652
rect 195244 50532 195296 50584
rect 368480 50532 368532 50584
rect 222384 50464 222436 50516
rect 462320 50464 462372 50516
rect 223764 50396 223816 50448
rect 465172 50396 465224 50448
rect 137284 50328 137336 50380
rect 178132 50328 178184 50380
rect 225052 50328 225104 50380
rect 473360 50328 473412 50380
rect 158904 49240 158956 49292
rect 258172 49240 258224 49292
rect 191288 49172 191340 49224
rect 354680 49172 354732 49224
rect 219624 49104 219676 49156
rect 451280 49104 451332 49156
rect 219532 49036 219584 49088
rect 455420 49036 455472 49088
rect 52460 48968 52512 49020
rect 95424 48968 95476 49020
rect 220912 48968 220964 49020
rect 458180 48968 458232 49020
rect 157616 47880 157668 47932
rect 253940 47880 253992 47932
rect 226984 47812 227036 47864
rect 440332 47812 440384 47864
rect 215300 47744 215352 47796
rect 440240 47744 440292 47796
rect 216772 47676 216824 47728
rect 444380 47676 444432 47728
rect 218244 47608 218296 47660
rect 448520 47608 448572 47660
rect 147956 47540 148008 47592
rect 219532 47540 219584 47592
rect 244464 47540 244516 47592
rect 535460 47540 535512 47592
rect 261484 46860 261536 46912
rect 550088 46860 550140 46912
rect 550548 46860 550600 46912
rect 157524 46452 157576 46504
rect 251456 46452 251508 46504
rect 192024 46384 192076 46436
rect 361580 46384 361632 46436
rect 196072 46316 196124 46368
rect 376760 46316 376812 46368
rect 204352 46248 204404 46300
rect 405740 46248 405792 46300
rect 207020 46180 207072 46232
rect 412640 46180 412692 46232
rect 550548 46180 550600 46232
rect 580172 46180 580224 46232
rect 169024 45092 169076 45144
rect 281540 45092 281592 45144
rect 189080 45024 189132 45076
rect 356060 45024 356112 45076
rect 193404 44956 193456 45008
rect 369860 44956 369912 45008
rect 138296 44888 138348 44940
rect 184204 44888 184256 44940
rect 211252 44888 211304 44940
rect 425060 44888 425112 44940
rect 30380 44820 30432 44872
rect 88524 44820 88576 44872
rect 145196 44820 145248 44872
rect 210516 44820 210568 44872
rect 229284 44820 229336 44872
rect 481640 44820 481692 44872
rect 156236 43732 156288 43784
rect 247040 43732 247092 43784
rect 211160 43664 211212 43716
rect 426440 43664 426492 43716
rect 73160 43596 73212 43648
rect 102324 43596 102376 43648
rect 215944 43596 215996 43648
rect 432052 43596 432104 43648
rect 66260 43528 66312 43580
rect 99564 43528 99616 43580
rect 212724 43528 212776 43580
rect 430580 43528 430632 43580
rect 59360 43460 59412 43512
rect 98276 43460 98328 43512
rect 214012 43460 214064 43512
rect 433340 43460 433392 43512
rect 22100 43392 22152 43444
rect 87236 43392 87288 43444
rect 102324 43392 102376 43444
rect 110696 43392 110748 43444
rect 145104 43392 145156 43444
rect 212632 43392 212684 43444
rect 236184 43392 236236 43444
rect 505100 43392 505152 43444
rect 171140 42304 171192 42356
rect 295340 42304 295392 42356
rect 193864 42236 193916 42288
rect 365720 42236 365772 42288
rect 35900 42168 35952 42220
rect 91192 42168 91244 42220
rect 208492 42168 208544 42220
rect 415400 42168 415452 42220
rect 16580 42100 16632 42152
rect 84384 42100 84436 42152
rect 209872 42100 209924 42152
rect 419540 42100 419592 42152
rect 1400 42032 1452 42084
rect 80336 42032 80388 42084
rect 125876 42032 125928 42084
rect 149152 42032 149204 42084
rect 149244 42032 149296 42084
rect 226524 42032 226576 42084
rect 229192 42032 229244 42084
rect 483020 42032 483072 42084
rect 162860 41012 162912 41064
rect 270500 41012 270552 41064
rect 167000 40944 167052 40996
rect 284392 40944 284444 40996
rect 94228 40876 94280 40928
rect 109132 40876 109184 40928
rect 202880 40876 202932 40928
rect 398932 40876 398984 40928
rect 129188 40808 129240 40860
rect 154856 40808 154908 40860
rect 216680 40808 216732 40860
rect 443000 40808 443052 40860
rect 44180 40740 44232 40792
rect 94136 40740 94188 40792
rect 135260 40740 135312 40792
rect 181076 40740 181128 40792
rect 242900 40740 242952 40792
rect 528560 40740 528612 40792
rect 20 40672 72 40724
rect 80244 40672 80296 40724
rect 145012 40672 145064 40724
rect 209872 40672 209924 40724
rect 252744 40672 252796 40724
rect 559012 40672 559064 40724
rect 198924 39584 198976 39636
rect 387800 39584 387852 39636
rect 200212 39516 200264 39568
rect 390560 39516 390612 39568
rect 206284 39448 206336 39500
rect 400220 39448 400272 39500
rect 204260 39380 204312 39432
rect 401600 39380 401652 39432
rect 154948 39312 155000 39364
rect 242900 39312 242952 39364
rect 244372 39312 244424 39364
rect 531412 39312 531464 39364
rect 153200 38224 153252 38276
rect 240324 38224 240376 38276
rect 194600 38156 194652 38208
rect 374092 38156 374144 38208
rect 197452 38088 197504 38140
rect 380900 38088 380952 38140
rect 198832 38020 198884 38072
rect 383660 38020 383712 38072
rect 217324 37952 217376 38004
rect 422300 37952 422352 38004
rect 237564 37884 237616 37936
rect 510620 37884 510672 37936
rect 152004 36864 152056 36916
rect 236184 36864 236236 36916
rect 186412 36796 186464 36848
rect 345020 36796 345072 36848
rect 191932 36728 191984 36780
rect 362960 36728 363012 36780
rect 193312 36660 193364 36712
rect 365812 36660 365864 36712
rect 214564 36592 214616 36644
rect 418160 36592 418212 36644
rect 236092 36524 236144 36576
rect 506572 36524 506624 36576
rect 191196 35436 191248 35488
rect 340880 35436 340932 35488
rect 183652 35368 183704 35420
rect 338120 35368 338172 35420
rect 140964 35300 141016 35352
rect 188436 35300 188488 35352
rect 254032 35300 254084 35352
rect 564624 35300 564676 35352
rect 147864 35232 147916 35284
rect 222384 35232 222436 35284
rect 256700 35232 256752 35284
rect 572812 35232 572864 35284
rect 151912 35164 151964 35216
rect 233424 35164 233476 35216
rect 256792 35164 256844 35216
rect 575480 35164 575532 35216
rect 180984 34008 181036 34060
rect 327080 34008 327132 34060
rect 182272 33940 182324 33992
rect 331220 33940 331272 33992
rect 182364 33872 182416 33924
rect 333980 33872 334032 33924
rect 213276 33804 213328 33856
rect 415492 33804 415544 33856
rect 147772 33736 147824 33788
rect 218244 33736 218296 33788
rect 226432 33736 226484 33788
rect 477500 33736 477552 33788
rect 176844 32648 176896 32700
rect 316040 32648 316092 32700
rect 178224 32580 178276 32632
rect 320180 32580 320232 32632
rect 179512 32512 179564 32564
rect 324412 32512 324464 32564
rect 213184 32444 213236 32496
rect 411260 32444 411312 32496
rect 146484 32376 146536 32428
rect 215300 32376 215352 32428
rect 218152 32376 218204 32428
rect 448612 32376 448664 32428
rect 173992 31288 174044 31340
rect 306380 31288 306432 31340
rect 175464 31220 175516 31272
rect 309140 31220 309192 31272
rect 176752 31152 176804 31204
rect 313280 31152 313332 31204
rect 139676 31084 139728 31136
rect 174544 31084 174596 31136
rect 209136 31084 209188 31136
rect 407120 31084 407172 31136
rect 143724 31016 143776 31068
rect 208492 31016 208544 31068
rect 224960 31016 225012 31068
rect 470600 31016 470652 31068
rect 165620 29928 165672 29980
rect 277400 29928 277452 29980
rect 172796 29860 172848 29912
rect 302240 29860 302292 29912
rect 195980 29792 196032 29844
rect 375380 29792 375432 29844
rect 138204 29724 138256 29776
rect 166356 29724 166408 29776
rect 251364 29724 251416 29776
rect 557540 29724 557592 29776
rect 142436 29656 142488 29708
rect 201592 29656 201644 29708
rect 252652 29656 252704 29708
rect 561864 29656 561916 29708
rect 142344 29588 142396 29640
rect 204260 29588 204312 29640
rect 255412 29588 255464 29640
rect 568580 29588 568632 29640
rect 161572 28568 161624 28620
rect 267832 28568 267884 28620
rect 164240 28500 164292 28552
rect 274640 28500 274692 28552
rect 192576 28432 192628 28484
rect 350540 28432 350592 28484
rect 244280 28364 244332 28416
rect 532700 28364 532752 28416
rect 136916 28296 136968 28348
rect 185032 28296 185084 28348
rect 249984 28296 250036 28348
rect 550640 28296 550692 28348
rect 140872 28228 140924 28280
rect 197452 28228 197504 28280
rect 251272 28228 251324 28280
rect 554780 28228 554832 28280
rect 160100 27208 160152 27260
rect 259644 27208 259696 27260
rect 161480 27140 161532 27192
rect 263600 27140 263652 27192
rect 197360 27072 197412 27124
rect 379520 27072 379572 27124
rect 132776 27004 132828 27056
rect 160744 27004 160796 27056
rect 237380 27004 237432 27056
rect 512000 27004 512052 27056
rect 139584 26936 139636 26988
rect 193312 26936 193364 26988
rect 241612 26936 241664 26988
rect 523132 26936 523184 26988
rect 150716 26868 150768 26920
rect 229192 26868 229244 26920
rect 241704 26868 241756 26920
rect 525800 26868 525852 26920
rect 156144 25848 156196 25900
rect 249984 25848 250036 25900
rect 157432 25780 157484 25832
rect 252652 25780 252704 25832
rect 186320 25712 186372 25764
rect 343640 25712 343692 25764
rect 233332 25644 233384 25696
rect 498292 25644 498344 25696
rect 234804 25576 234856 25628
rect 500960 25576 501012 25628
rect 138112 25508 138164 25560
rect 190644 25508 190696 25560
rect 236000 25508 236052 25560
rect 507860 25508 507912 25560
rect 154764 24488 154816 24540
rect 242992 24488 243044 24540
rect 156052 24420 156104 24472
rect 245844 24420 245896 24472
rect 212540 24352 212592 24404
rect 429200 24352 429252 24404
rect 230664 24284 230716 24336
rect 487160 24284 487212 24336
rect 230756 24216 230808 24268
rect 489920 24216 489972 24268
rect 134524 24148 134576 24200
rect 167000 24148 167052 24200
rect 231952 24148 232004 24200
rect 494060 24148 494112 24200
rect 136824 24080 136876 24132
rect 183652 24080 183704 24132
rect 241520 24080 241572 24132
rect 524420 24080 524472 24132
rect 110696 23400 110748 23452
rect 113364 23400 113416 23452
rect 158812 22924 158864 22976
rect 256700 22924 256752 22976
rect 218060 22856 218112 22908
rect 449900 22856 449952 22908
rect 227812 22788 227864 22840
rect 480260 22788 480312 22840
rect 53840 22720 53892 22772
rect 96804 22720 96856 22772
rect 141424 22720 141476 22772
rect 168472 22720 168524 22772
rect 240232 22720 240284 22772
rect 521660 22720 521712 22772
rect 103888 22108 103940 22160
rect 112076 22108 112128 22160
rect 178040 21632 178092 21684
rect 318800 21632 318852 21684
rect 182180 21564 182232 21616
rect 332692 21564 332744 21616
rect 144184 21496 144236 21548
rect 179512 21496 179564 21548
rect 183560 21496 183612 21548
rect 336740 21496 336792 21548
rect 132684 21428 132736 21480
rect 172796 21428 172848 21480
rect 184940 21428 184992 21480
rect 340972 21428 341024 21480
rect 77300 21360 77352 21412
rect 103796 21360 103848 21412
rect 134064 21360 134116 21412
rect 176752 21360 176804 21412
rect 210424 21360 210476 21412
rect 404360 21360 404412 21412
rect 3424 20612 3476 20664
rect 560116 20612 560168 20664
rect 560944 20612 560996 20664
rect 579988 20612 580040 20664
rect 172704 20204 172756 20256
rect 300860 20204 300912 20256
rect 173900 20136 173952 20188
rect 305000 20136 305052 20188
rect 133972 20068 134024 20120
rect 162124 20068 162176 20120
rect 175280 20068 175332 20120
rect 307852 20068 307904 20120
rect 132592 20000 132644 20052
rect 160836 20000 160888 20052
rect 175372 20000 175424 20052
rect 311900 20000 311952 20052
rect 98276 19932 98328 19984
rect 110604 19932 110656 19984
rect 130016 19932 130068 19984
rect 161480 19932 161532 19984
rect 207664 19932 207716 19984
rect 397460 19932 397512 19984
rect 179420 18844 179472 18896
rect 322940 18844 322992 18896
rect 188344 18776 188396 18828
rect 238760 18776 238812 18828
rect 245752 18776 245804 18828
rect 539692 18776 539744 18828
rect 144920 18708 144972 18760
rect 214012 18708 214064 18760
rect 252560 18708 252612 18760
rect 560300 18708 560352 18760
rect 150624 18640 150676 18692
rect 231952 18640 232004 18692
rect 255320 18640 255372 18692
rect 567200 18640 567252 18692
rect 24860 18572 24912 18624
rect 87144 18572 87196 18624
rect 124496 18572 124548 18624
rect 144920 18572 144972 18624
rect 151820 18572 151872 18624
rect 234804 18572 234856 18624
rect 258080 18572 258132 18624
rect 578240 18572 578292 18624
rect 180892 17484 180944 17536
rect 325700 17484 325752 17536
rect 60740 17416 60792 17468
rect 98184 17416 98236 17468
rect 123024 17416 123076 17468
rect 142344 17416 142396 17468
rect 231860 17416 231912 17468
rect 492680 17416 492732 17468
rect 45560 17348 45612 17400
rect 94044 17348 94096 17400
rect 139492 17348 139544 17400
rect 195980 17348 196032 17400
rect 233240 17348 233292 17400
rect 496820 17348 496872 17400
rect 38660 17280 38712 17332
rect 91284 17280 91336 17332
rect 140780 17280 140832 17332
rect 200212 17280 200264 17332
rect 234712 17280 234764 17332
rect 499580 17280 499632 17332
rect 15200 17212 15252 17264
rect 84292 17212 84344 17264
rect 142252 17212 142304 17264
rect 202880 17212 202932 17264
rect 234620 17212 234672 17264
rect 503720 17212 503772 17264
rect 191104 16124 191156 16176
rect 348056 16124 348108 16176
rect 75000 16056 75052 16108
rect 100024 16056 100076 16108
rect 166264 16056 166316 16108
rect 182180 16056 182232 16108
rect 205732 16056 205784 16108
rect 407212 16056 407264 16108
rect 67640 15988 67692 16040
rect 100944 15988 100996 16040
rect 136732 15988 136784 16040
rect 170404 15988 170456 16040
rect 205824 15988 205876 16040
rect 410800 15988 410852 16040
rect 31944 15920 31996 15972
rect 89904 15920 89956 15972
rect 133880 15920 133932 15972
rect 175464 15920 175516 15972
rect 208400 15920 208452 15972
rect 417424 15920 417476 15972
rect 24216 15852 24268 15904
rect 87052 15852 87104 15904
rect 122932 15852 122984 15904
rect 138848 15852 138900 15904
rect 139400 15852 139452 15904
rect 193404 15852 193456 15904
rect 223580 15852 223632 15904
rect 467472 15852 467524 15904
rect 190552 14696 190604 14748
rect 361120 14696 361172 14748
rect 56784 14628 56836 14680
rect 96712 14628 96764 14680
rect 191840 14628 191892 14680
rect 364616 14628 364668 14680
rect 53012 14560 53064 14612
rect 93124 14560 93176 14612
rect 129832 14560 129884 14612
rect 160652 14560 160704 14612
rect 193220 14560 193272 14612
rect 367744 14560 367796 14612
rect 14280 14492 14332 14544
rect 84200 14492 84252 14544
rect 129924 14492 129976 14544
rect 164424 14492 164476 14544
rect 200120 14492 200172 14544
rect 390652 14492 390704 14544
rect 9680 14424 9732 14476
rect 83004 14424 83056 14476
rect 85764 14424 85816 14476
rect 101404 14424 101456 14476
rect 132500 14424 132552 14476
rect 171968 14424 172020 14476
rect 222292 14424 222344 14476
rect 463976 14424 464028 14476
rect 157340 13404 157392 13456
rect 251272 13404 251324 13456
rect 172612 13336 172664 13388
rect 299480 13336 299532 13388
rect 69848 13268 69900 13320
rect 100852 13268 100904 13320
rect 158720 13268 158772 13320
rect 255872 13268 255924 13320
rect 255964 13268 256016 13320
rect 454040 13268 454092 13320
rect 41880 13200 41932 13252
rect 92664 13200 92716 13252
rect 128360 13200 128412 13252
rect 157800 13200 157852 13252
rect 222200 13200 222252 13252
rect 459928 13200 459980 13252
rect 34520 13132 34572 13184
rect 89812 13132 89864 13184
rect 128452 13132 128504 13184
rect 158904 13132 158956 13184
rect 226340 13132 226392 13184
rect 474096 13132 474148 13184
rect 27712 13064 27764 13116
rect 88432 13064 88484 13116
rect 118884 13064 118936 13116
rect 128176 13064 128228 13116
rect 129740 13064 129792 13116
rect 163688 13064 163740 13116
rect 249892 13064 249944 13116
rect 550272 13064 550324 13116
rect 143540 12724 143592 12776
rect 143724 12724 143776 12776
rect 234804 12724 234856 12776
rect 235816 12724 235868 12776
rect 176660 11976 176712 12028
rect 316224 11976 316276 12028
rect 61568 11908 61620 11960
rect 98092 11908 98144 11960
rect 230572 11908 230624 11960
rect 490012 11908 490064 11960
rect 63224 11840 63276 11892
rect 99472 11840 99524 11892
rect 125784 11840 125836 11892
rect 150624 11840 150676 11892
rect 154672 11840 154724 11892
rect 241704 11840 241756 11892
rect 44272 11772 44324 11824
rect 92572 11772 92624 11824
rect 127164 11772 127216 11824
rect 153752 11772 153804 11824
rect 154580 11772 154632 11824
rect 245200 11840 245252 11892
rect 248512 11840 248564 11892
rect 548616 11840 548668 11892
rect 242900 11772 242952 11824
rect 244096 11772 244148 11824
rect 249800 11772 249852 11824
rect 552664 11772 552716 11824
rect 17960 11704 18012 11756
rect 85672 11704 85724 11756
rect 89168 11704 89220 11756
rect 105544 11704 105596 11756
rect 125692 11704 125744 11756
rect 151820 11704 151872 11756
rect 155960 11704 156012 11756
rect 248512 11704 248564 11756
rect 251180 11704 251232 11756
rect 556252 11704 556304 11756
rect 117412 10956 117464 11008
rect 120632 10956 120684 11008
rect 150532 10616 150584 10668
rect 231032 10616 231084 10668
rect 192484 10548 192536 10600
rect 357532 10548 357584 10600
rect 56048 10480 56100 10532
rect 96620 10480 96672 10532
rect 220820 10480 220872 10532
rect 456892 10480 456944 10532
rect 40224 10412 40276 10464
rect 92756 10412 92808 10464
rect 129096 10412 129148 10464
rect 143540 10412 143592 10464
rect 227720 10412 227772 10464
rect 481732 10412 481784 10464
rect 13544 10344 13596 10396
rect 82912 10344 82964 10396
rect 92572 10344 92624 10396
rect 107016 10344 107068 10396
rect 122840 10344 122892 10396
rect 141240 10344 141292 10396
rect 146392 10344 146444 10396
rect 216864 10344 216916 10396
rect 229100 10344 229152 10396
rect 484768 10344 484820 10396
rect 3608 10276 3660 10328
rect 80152 10276 80204 10328
rect 87512 10276 87564 10328
rect 106372 10276 106424 10328
rect 125600 10276 125652 10328
rect 147864 10276 147916 10328
rect 149060 10276 149112 10328
rect 227536 10276 227588 10328
rect 230480 10276 230532 10328
rect 488816 10276 488868 10328
rect 116216 9596 116268 9648
rect 118792 9596 118844 9648
rect 143632 9256 143684 9308
rect 209780 9256 209832 9308
rect 86868 9188 86920 9240
rect 106464 9188 106516 9240
rect 198740 9188 198792 9240
rect 387156 9188 387208 9240
rect 72608 9120 72660 9172
rect 102232 9120 102284 9172
rect 118884 9120 118936 9172
rect 129372 9120 129424 9172
rect 201500 9120 201552 9172
rect 395344 9120 395396 9172
rect 58440 9052 58492 9104
rect 98000 9052 98052 9104
rect 124404 9052 124456 9104
rect 144736 9052 144788 9104
rect 205640 9052 205692 9104
rect 409604 9052 409656 9104
rect 30104 8984 30156 9036
rect 88616 8984 88668 9036
rect 123484 8984 123536 9036
rect 134156 8984 134208 9036
rect 142160 8984 142212 9036
rect 202696 8984 202748 9036
rect 209872 8984 209924 9036
rect 423772 8984 423824 9036
rect 26516 8916 26568 8968
rect 86960 8916 87012 8968
rect 101036 8916 101088 8968
rect 110512 8916 110564 8968
rect 122104 8916 122156 8968
rect 132960 8916 133012 8968
rect 143724 8916 143776 8968
rect 206192 8916 206244 8968
rect 219440 8916 219492 8968
rect 453304 8916 453356 8968
rect 117320 8236 117372 8288
rect 122288 8236 122340 8288
rect 82084 7828 82136 7880
rect 97264 7828 97316 7880
rect 187700 7828 187752 7880
rect 349252 7828 349304 7880
rect 47860 7760 47912 7812
rect 93952 7760 94004 7812
rect 121552 7760 121604 7812
rect 137652 7760 137704 7812
rect 187792 7760 187844 7812
rect 352840 7760 352892 7812
rect 21824 7692 21876 7744
rect 85856 7692 85908 7744
rect 97448 7692 97500 7744
rect 109224 7692 109276 7744
rect 138020 7692 138072 7744
rect 188528 7692 188580 7744
rect 190460 7692 190512 7744
rect 359924 7692 359976 7744
rect 7656 7624 7708 7676
rect 81624 7624 81676 7676
rect 90364 7624 90416 7676
rect 107844 7624 107896 7676
rect 121644 7624 121696 7676
rect 135260 7624 135312 7676
rect 136640 7624 136692 7676
rect 187332 7624 187384 7676
rect 209044 7624 209096 7676
rect 394240 7624 394292 7676
rect 2872 7556 2924 7608
rect 80060 7556 80112 7608
rect 80888 7556 80940 7608
rect 105084 7556 105136 7608
rect 130568 7556 130620 7608
rect 561680 7556 561732 7608
rect 561312 6808 561364 6860
rect 580172 6808 580224 6860
rect 169760 6400 169812 6452
rect 292580 6400 292632 6452
rect 77392 6332 77444 6384
rect 103704 6332 103756 6384
rect 131212 6332 131264 6384
rect 169576 6332 169628 6384
rect 172520 6332 172572 6384
rect 299664 6332 299716 6384
rect 48964 6264 49016 6316
rect 93860 6264 93912 6316
rect 126980 6264 127032 6316
rect 127164 6264 127216 6316
rect 203524 6264 203576 6316
rect 383568 6264 383620 6316
rect 33600 6196 33652 6248
rect 89720 6196 89772 6248
rect 91560 6196 91612 6248
rect 107752 6196 107804 6248
rect 131120 6196 131172 6248
rect 166080 6196 166132 6248
rect 168380 6196 168432 6248
rect 288992 6196 289044 6248
rect 289084 6196 289136 6248
rect 475752 6196 475804 6248
rect 8760 6128 8812 6180
rect 81532 6128 81584 6180
rect 84476 6128 84528 6180
rect 104992 6128 105044 6180
rect 126980 6128 127032 6180
rect 561772 6128 561824 6180
rect 127072 5924 127124 5976
rect 128360 5924 128412 5976
rect 126244 5516 126296 5568
rect 131764 5516 131816 5568
rect 83280 5108 83332 5160
rect 105176 5108 105228 5160
rect 187056 5108 187108 5160
rect 225144 5108 225196 5160
rect 79692 5040 79744 5092
rect 103612 5040 103664 5092
rect 180800 5040 180852 5092
rect 330392 5040 330444 5092
rect 76196 4972 76248 5024
rect 103520 4972 103572 5024
rect 213920 4972 213972 5024
rect 437940 4972 437992 5024
rect 69112 4904 69164 4956
rect 100944 4904 100996 4956
rect 118700 4904 118752 4956
rect 125876 4904 125928 4956
rect 129004 4904 129056 4956
rect 140044 4904 140096 4956
rect 146300 4904 146352 4956
rect 218060 4904 218112 4956
rect 240140 4904 240192 4956
rect 519544 4972 519596 5024
rect 65616 4836 65668 4888
rect 99656 4836 99708 4888
rect 121460 4836 121512 4888
rect 136456 4836 136508 4888
rect 147680 4836 147732 4888
rect 221556 4836 221608 4888
rect 245660 4836 245712 4888
rect 537208 4836 537260 4888
rect 12348 4768 12400 4820
rect 83096 4768 83148 4820
rect 124312 4768 124364 4820
rect 147128 4768 147180 4820
rect 150440 4768 150492 4820
rect 228732 4768 228784 4820
rect 248420 4768 248472 4820
rect 547880 4768 547932 4820
rect 105728 4156 105780 4208
rect 111984 4156 112036 4208
rect 64328 4088 64380 4140
rect 65524 4088 65576 4140
rect 119344 4088 119396 4140
rect 123484 4088 123536 4140
rect 170404 3748 170456 3800
rect 162124 3680 162176 3732
rect 20628 3612 20680 3664
rect 28264 3612 28316 3664
rect 11152 3544 11204 3596
rect 15844 3544 15896 3596
rect 43076 3544 43128 3596
rect 53104 3544 53156 3596
rect 99840 3544 99892 3596
rect 109684 3612 109736 3664
rect 160744 3612 160796 3664
rect 5264 3476 5316 3528
rect 10324 3476 10376 3528
rect 28908 3476 28960 3528
rect 32404 3476 32456 3528
rect 44180 3476 44232 3528
rect 45100 3476 45152 3528
rect 6460 3408 6512 3460
rect 35992 3340 36044 3392
rect 50344 3476 50396 3528
rect 102140 3476 102192 3528
rect 103336 3476 103388 3528
rect 103428 3476 103480 3528
rect 108304 3544 108356 3596
rect 109316 3544 109368 3596
rect 111064 3544 111116 3596
rect 128360 3544 128412 3596
rect 153016 3544 153068 3596
rect 160836 3544 160888 3596
rect 170772 3544 170824 3596
rect 407764 3748 407816 3800
rect 461584 3748 461636 3800
rect 188436 3680 188488 3732
rect 199108 3680 199160 3732
rect 411996 3680 412048 3732
rect 468668 3680 468720 3732
rect 186136 3612 186188 3664
rect 193312 3612 193364 3664
rect 194416 3612 194468 3664
rect 258724 3612 258776 3664
rect 177856 3544 177908 3596
rect 186964 3544 187016 3596
rect 207388 3544 207440 3596
rect 210516 3544 210568 3596
rect 212172 3544 212224 3596
rect 251272 3544 251324 3596
rect 252376 3544 252428 3596
rect 259460 3544 259512 3596
rect 106924 3476 106976 3528
rect 111892 3476 111944 3528
rect 116124 3476 116176 3528
rect 117596 3476 117648 3528
rect 135904 3476 135956 3528
rect 160100 3476 160152 3528
rect 174268 3476 174320 3528
rect 174544 3476 174596 3528
rect 195612 3476 195664 3528
rect 81808 3408 81860 3460
rect 93952 3340 94004 3392
rect 106832 3408 106884 3460
rect 116032 3408 116084 3460
rect 119896 3408 119948 3460
rect 127164 3408 127216 3460
rect 156604 3408 156656 3460
rect 166356 3408 166408 3460
rect 192024 3408 192076 3460
rect 422944 3612 422996 3664
rect 583392 3612 583444 3664
rect 267740 3544 267792 3596
rect 268476 3544 268528 3596
rect 276020 3544 276072 3596
rect 276756 3544 276808 3596
rect 307852 3544 307904 3596
rect 309048 3544 309100 3596
rect 316040 3544 316092 3596
rect 317328 3544 317380 3596
rect 324320 3544 324372 3596
rect 325608 3544 325660 3596
rect 332692 3544 332744 3596
rect 333888 3544 333940 3596
rect 357532 3544 357584 3596
rect 358728 3544 358780 3596
rect 365812 3544 365864 3596
rect 367008 3544 367060 3596
rect 374000 3544 374052 3596
rect 375288 3544 375340 3596
rect 390560 3544 390612 3596
rect 391848 3544 391900 3596
rect 398840 3544 398892 3596
rect 400128 3544 400180 3596
rect 418804 3544 418856 3596
rect 581000 3544 581052 3596
rect 479340 3476 479392 3528
rect 481640 3476 481692 3528
rect 482468 3476 482520 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 498200 3476 498252 3528
rect 499028 3476 499080 3528
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 523040 3476 523092 3528
rect 523868 3476 523920 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 556160 3476 556212 3528
rect 556988 3476 557040 3528
rect 572720 3476 572772 3528
rect 573548 3476 573600 3528
rect 582196 3408 582248 3460
rect 423680 3340 423732 3392
rect 424968 3340 425020 3392
rect 432052 3340 432104 3392
rect 433248 3340 433300 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 96252 3272 96304 3324
rect 103428 3272 103480 3324
rect 19432 3000 19484 3052
rect 25504 3000 25556 3052
rect 184204 2932 184256 2984
rect 189724 2932 189776 2984
rect 415400 2864 415452 2916
rect 416688 2864 416740 2916
rect 299480 2728 299532 2780
rect 300768 2728 300820 2780
rect 407120 2592 407172 2644
rect 408408 2592 408460 2644
rect 340880 2320 340932 2372
rect 342168 2320 342220 2372
rect 349160 2320 349212 2372
rect 350448 2320 350500 2372
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3436 424386 3464 632023
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3514 475688 3570 475697
rect 3514 475623 3570 475632
rect 3528 425814 3556 475623
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3620 428466 3648 462567
rect 3698 449576 3754 449585
rect 3698 449511 3754 449520
rect 3608 428460 3660 428466
rect 3608 428402 3660 428408
rect 3712 427106 3740 449511
rect 3700 427100 3752 427106
rect 3700 427042 3752 427048
rect 3516 425808 3568 425814
rect 3516 425750 3568 425756
rect 3424 424380 3476 424386
rect 3424 424322 3476 424328
rect 4896 423700 4948 423706
rect 4896 423642 4948 423648
rect 4066 423600 4122 423609
rect 4066 423535 4122 423544
rect 4080 423026 4108 423535
rect 4802 423192 4858 423201
rect 4802 423127 4858 423136
rect 4068 423020 4120 423026
rect 4068 422962 4120 422968
rect 3514 422512 3570 422521
rect 3514 422447 3570 422456
rect 3422 421696 3478 421705
rect 3422 421631 3478 421640
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3056 358760 3108 358766
rect 3056 358702 3108 358708
rect 3068 358465 3096 358702
rect 3054 358456 3110 358465
rect 3054 358391 3110 358400
rect 2964 346384 3016 346390
rect 2964 346326 3016 346332
rect 2976 345409 3004 346326
rect 2962 345400 3018 345409
rect 2962 345335 3018 345344
rect 3332 319456 3384 319462
rect 3332 319398 3384 319404
rect 3344 319297 3372 319398
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3240 293956 3292 293962
rect 3240 293898 3292 293904
rect 3252 293185 3280 293898
rect 3238 293176 3294 293185
rect 3238 293111 3294 293120
rect 3330 267200 3386 267209
rect 3330 267135 3386 267144
rect 3344 267034 3372 267135
rect 3332 267028 3384 267034
rect 3332 266970 3384 266976
rect 2964 255264 3016 255270
rect 2964 255206 3016 255212
rect 2976 254153 3004 255206
rect 2962 254144 3018 254153
rect 2962 254079 3018 254088
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 214606 3372 214911
rect 3332 214600 3384 214606
rect 3332 214542 3384 214548
rect 2780 162988 2832 162994
rect 2780 162930 2832 162936
rect 2792 162897 2820 162930
rect 2778 162888 2834 162897
rect 2778 162823 2834 162832
rect 2780 150204 2832 150210
rect 2780 150146 2832 150152
rect 2792 149841 2820 150146
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 2964 85536 3016 85542
rect 2964 85478 3016 85484
rect 2976 84697 3004 85478
rect 2962 84688 3018 84697
rect 2962 84623 3018 84632
rect 3436 45529 3464 421631
rect 3528 188873 3556 422447
rect 3606 421832 3662 421841
rect 3606 421767 3662 421776
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3620 58585 3648 421767
rect 3700 421660 3752 421666
rect 3700 421602 3752 421608
rect 3712 201929 3740 421602
rect 3884 421592 3936 421598
rect 3790 421560 3846 421569
rect 3884 421534 3936 421540
rect 3790 421495 3846 421504
rect 3804 241097 3832 421495
rect 3896 397497 3924 421534
rect 3882 397488 3938 397497
rect 3882 397423 3938 397432
rect 3790 241088 3846 241097
rect 3790 241023 3846 241032
rect 3698 201920 3754 201929
rect 3698 201855 3754 201864
rect 3792 201544 3844 201550
rect 3792 201486 3844 201492
rect 3700 200320 3752 200326
rect 3700 200262 3752 200268
rect 3712 71641 3740 200262
rect 3698 71632 3754 71641
rect 3698 71567 3754 71576
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 1400 42084 1452 42090
rect 1400 42026 1452 42032
rect 20 40724 72 40730
rect 20 40666 72 40672
rect 32 16574 60 40666
rect 32 16546 152 16574
rect 124 354 152 16546
rect 542 354 654 480
rect 124 326 654 354
rect 1412 354 1440 42026
rect 3804 32473 3832 201486
rect 3884 200388 3936 200394
rect 3884 200330 3936 200336
rect 3896 110673 3924 200330
rect 3882 110664 3938 110673
rect 3882 110599 3938 110608
rect 4816 97782 4844 423127
rect 4908 423026 4936 423642
rect 4896 423020 4948 423026
rect 4896 422962 4948 422968
rect 4908 203590 4936 422962
rect 4986 422648 5042 422657
rect 4986 422583 5042 422592
rect 4896 203584 4948 203590
rect 4896 203526 4948 203532
rect 4896 200456 4948 200462
rect 4896 200398 4948 200404
rect 4908 162994 4936 200398
rect 4896 162988 4948 162994
rect 4896 162930 4948 162936
rect 5000 150210 5028 422583
rect 40052 203726 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 427174 71820 702986
rect 89180 700466 89208 703520
rect 105464 700534 105492 703520
rect 105452 700528 105504 700534
rect 105452 700470 105504 700476
rect 89168 700460 89220 700466
rect 89168 700402 89220 700408
rect 71780 427168 71832 427174
rect 71780 427110 71832 427116
rect 136652 425746 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 153212 599622 153240 702406
rect 170324 700602 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 170312 700596 170364 700602
rect 170312 700538 170364 700544
rect 180064 700596 180116 700602
rect 180064 700538 180116 700544
rect 153200 599616 153252 599622
rect 153200 599558 153252 599564
rect 177304 565888 177356 565894
rect 177304 565830 177356 565836
rect 177316 428534 177344 565830
rect 177396 514820 177448 514826
rect 177396 514762 177448 514768
rect 177408 428602 177436 514762
rect 177396 428596 177448 428602
rect 177396 428538 177448 428544
rect 177304 428528 177356 428534
rect 177304 428470 177356 428476
rect 136640 425740 136692 425746
rect 136640 425682 136692 425688
rect 180076 423842 180104 700538
rect 185584 700528 185636 700534
rect 185584 700470 185636 700476
rect 185596 425610 185624 700470
rect 193864 683188 193916 683194
rect 193864 683130 193916 683136
rect 184940 425604 184992 425610
rect 184940 425546 184992 425552
rect 185584 425604 185636 425610
rect 185584 425546 185636 425552
rect 179420 423836 179472 423842
rect 179420 423778 179472 423784
rect 180064 423836 180116 423842
rect 180064 423778 180116 423784
rect 77944 423768 77996 423774
rect 77944 423710 77996 423716
rect 43444 422952 43496 422958
rect 43444 422894 43496 422900
rect 43456 411262 43484 422894
rect 43444 411256 43496 411262
rect 43444 411198 43496 411204
rect 40040 203720 40092 203726
rect 40040 203662 40092 203668
rect 4988 150204 5040 150210
rect 4988 150146 5040 150152
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 77956 85542 77984 423710
rect 175924 423088 175976 423094
rect 175924 423030 175976 423036
rect 87604 423020 87656 423026
rect 87604 422962 87656 422968
rect 79322 422784 79378 422793
rect 79322 422719 79378 422728
rect 79336 137970 79364 422719
rect 87616 358766 87644 422962
rect 126980 422000 127032 422006
rect 126980 421942 127032 421948
rect 87604 358760 87656 358766
rect 87604 358702 87656 358708
rect 113180 298784 113232 298790
rect 113180 298726 113232 298732
rect 109040 224256 109092 224262
rect 109040 224198 109092 224204
rect 103980 206304 104032 206310
rect 103980 206246 104032 206252
rect 100024 201680 100076 201686
rect 100024 201622 100076 201628
rect 95148 201612 95200 201618
rect 95148 201554 95200 201560
rect 85488 200524 85540 200530
rect 85488 200466 85540 200472
rect 81072 200184 81124 200190
rect 81072 200126 81124 200132
rect 81084 199866 81112 200126
rect 85500 199866 85528 200466
rect 90548 200252 90600 200258
rect 90548 200194 90600 200200
rect 90560 199866 90588 200194
rect 95160 199866 95188 201554
rect 100036 199866 100064 201622
rect 80776 199838 81112 199866
rect 85468 199838 85528 199866
rect 90252 199838 90588 199866
rect 94944 199838 95188 199866
rect 99728 199838 100064 199866
rect 103992 199866 104020 206246
rect 109052 199866 109080 224198
rect 113192 209774 113220 298726
rect 126992 209774 127020 421942
rect 136640 421728 136692 421734
rect 136640 421670 136692 421676
rect 132500 420164 132552 420170
rect 132500 420106 132552 420112
rect 113192 209746 113496 209774
rect 126992 209746 127756 209774
rect 113468 199866 113496 209746
rect 123668 202564 123720 202570
rect 123668 202506 123720 202512
rect 118976 202156 119028 202162
rect 118976 202098 119028 202104
rect 118988 199866 119016 202098
rect 123680 199866 123708 202506
rect 103992 199838 104420 199866
rect 109052 199838 109204 199866
rect 113468 199838 113896 199866
rect 118680 199838 119016 199866
rect 123372 199838 123708 199866
rect 127728 199866 127756 209746
rect 132512 199866 132540 420106
rect 136652 209774 136680 421670
rect 160100 420096 160152 420102
rect 160100 420038 160152 420044
rect 160112 209774 160140 420038
rect 175936 306338 175964 423030
rect 175924 306332 175976 306338
rect 175924 306274 175976 306280
rect 179432 209774 179460 423778
rect 184952 209774 184980 425546
rect 185596 425134 185624 425546
rect 185584 425128 185636 425134
rect 185584 425070 185636 425076
rect 193876 419694 193904 683130
rect 201512 427242 201540 702986
rect 218992 699718 219020 703520
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 220084 699712 220136 699718
rect 220084 699654 220136 699660
rect 202880 579692 202932 579698
rect 202880 579634 202932 579640
rect 201500 427236 201552 427242
rect 201500 427178 201552 427184
rect 198740 424380 198792 424386
rect 198740 424322 198792 424328
rect 198752 423910 198780 424322
rect 198740 423904 198792 423910
rect 198740 423846 198792 423852
rect 193864 419688 193916 419694
rect 193864 419630 193916 419636
rect 193876 419558 193904 419630
rect 193220 419552 193272 419558
rect 193220 419494 193272 419500
rect 193864 419552 193916 419558
rect 193864 419494 193916 419500
rect 193232 209774 193260 419494
rect 136652 209746 137232 209774
rect 160112 209746 160876 209774
rect 179432 209746 179828 209774
rect 184952 209746 185072 209774
rect 193232 209746 194088 209774
rect 137204 199866 137232 209746
rect 156880 202496 156932 202502
rect 156880 202438 156932 202444
rect 152096 202428 152148 202434
rect 152096 202370 152148 202376
rect 147404 202360 147456 202366
rect 147404 202302 147456 202308
rect 142620 202292 142672 202298
rect 142620 202234 142672 202240
rect 142632 199866 142660 202234
rect 147416 199866 147444 202302
rect 152108 199866 152136 202370
rect 156892 199866 156920 202438
rect 127728 199838 128156 199866
rect 132512 199838 132848 199866
rect 137204 199838 137632 199866
rect 142324 199838 142660 199866
rect 147108 199838 147444 199866
rect 151800 199838 152136 199866
rect 156584 199838 156920 199866
rect 160848 199866 160876 209746
rect 170312 203788 170364 203794
rect 170312 203730 170364 203736
rect 165620 203652 165672 203658
rect 165620 203594 165672 203600
rect 165632 199866 165660 203594
rect 170324 199866 170352 203730
rect 175832 202224 175884 202230
rect 175832 202166 175884 202172
rect 175844 199866 175872 202166
rect 160848 199838 161276 199866
rect 165632 199838 166060 199866
rect 170324 199838 170752 199866
rect 175536 199838 175872 199866
rect 179800 199866 179828 209746
rect 179800 199838 180228 199866
rect 185044 199730 185072 209746
rect 189080 203720 189132 203726
rect 189080 203662 189132 203668
rect 189092 202842 189120 203662
rect 189080 202836 189132 202842
rect 189080 202778 189132 202784
rect 189724 202836 189776 202842
rect 189724 202778 189776 202784
rect 189736 199866 189764 202778
rect 189704 199838 189764 199866
rect 194060 199866 194088 209746
rect 198752 199866 198780 423846
rect 202892 209774 202920 579634
rect 208400 527196 208452 527202
rect 208400 527138 208452 527144
rect 202892 209746 203564 209774
rect 203536 199866 203564 209746
rect 208412 199866 208440 527138
rect 220096 428670 220124 699654
rect 220084 428664 220136 428670
rect 220084 428606 220136 428612
rect 212540 425808 212592 425814
rect 212540 425750 212592 425756
rect 212552 425202 212580 425750
rect 212540 425196 212592 425202
rect 212540 425138 212592 425144
rect 212552 209774 212580 425138
rect 234632 425066 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 266372 425814 266400 697546
rect 282932 497486 282960 702406
rect 299492 511970 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 299480 511964 299532 511970
rect 299480 511906 299532 511912
rect 300124 511964 300176 511970
rect 300124 511906 300176 511912
rect 300136 510678 300164 511906
rect 300124 510672 300176 510678
rect 300124 510614 300176 510620
rect 282920 497480 282972 497486
rect 282920 497422 282972 497428
rect 266360 425808 266412 425814
rect 266360 425750 266412 425756
rect 234620 425060 234672 425066
rect 234620 425002 234672 425008
rect 235264 425060 235316 425066
rect 235264 425002 235316 425008
rect 235276 423978 235304 425002
rect 235264 423972 235316 423978
rect 235264 423914 235316 423920
rect 232504 420232 232556 420238
rect 232504 420174 232556 420180
rect 226982 419928 227038 419937
rect 226982 419863 227038 419872
rect 222200 371272 222252 371278
rect 223488 371272 223540 371278
rect 222200 371214 222252 371220
rect 223486 371240 223488 371249
rect 223540 371240 223542 371249
rect 222212 209774 222240 371214
rect 223486 371175 223542 371184
rect 226996 320142 227024 419863
rect 226340 320136 226392 320142
rect 226340 320078 226392 320084
rect 226984 320136 227036 320142
rect 226984 320078 227036 320084
rect 226352 319462 226380 320078
rect 226340 319456 226392 319462
rect 226340 319398 226392 319404
rect 226352 209774 226380 319398
rect 232516 267238 232544 420174
rect 231860 267232 231912 267238
rect 231860 267174 231912 267180
rect 232504 267232 232556 267238
rect 232504 267174 232556 267180
rect 231872 267034 231900 267174
rect 231860 267028 231912 267034
rect 231860 266970 231912 266976
rect 231872 209774 231900 266970
rect 212552 209746 213040 209774
rect 222212 209746 222516 209774
rect 226352 209746 227208 209774
rect 231872 209746 231992 209774
rect 213012 199866 213040 209746
rect 218152 203584 218204 203590
rect 218152 203526 218204 203532
rect 194060 199838 194488 199866
rect 198752 199838 199180 199866
rect 203536 199838 203964 199866
rect 208412 199838 208656 199866
rect 213012 199838 213440 199866
rect 218164 199730 218192 203526
rect 222488 199866 222516 209746
rect 227180 199866 227208 209746
rect 231964 199866 231992 209746
rect 235276 202230 235304 423914
rect 284944 421932 284996 421938
rect 284944 421874 284996 421880
rect 236644 419756 236696 419762
rect 236644 419698 236696 419704
rect 236656 214606 236684 419698
rect 236000 214600 236052 214606
rect 236000 214542 236052 214548
rect 236644 214600 236696 214606
rect 236644 214542 236696 214548
rect 236012 209774 236040 214542
rect 236012 209746 236684 209774
rect 235264 202224 235316 202230
rect 235264 202166 235316 202172
rect 236656 199866 236684 209746
rect 284956 202570 284984 421874
rect 300136 203794 300164 510614
rect 331232 425882 331260 702986
rect 348804 700126 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700120 348844 700126
rect 348792 700062 348844 700068
rect 349804 700120 349856 700126
rect 349804 700062 349856 700068
rect 349816 428738 349844 700062
rect 349804 428732 349856 428738
rect 349804 428674 349856 428680
rect 364352 426426 364380 702406
rect 397472 427310 397500 703520
rect 412652 428806 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 412640 428800 412692 428806
rect 412640 428742 412692 428748
rect 397460 427304 397512 427310
rect 397460 427246 397512 427252
rect 364340 426420 364392 426426
rect 364340 426362 364392 426368
rect 364984 426420 365036 426426
rect 364984 426362 365036 426368
rect 331220 425876 331272 425882
rect 331220 425818 331272 425824
rect 364996 425270 365024 426362
rect 364984 425264 365036 425270
rect 364984 425206 365036 425212
rect 352564 422544 352616 422550
rect 352564 422486 352616 422492
rect 352576 255270 352604 422486
rect 352564 255264 352616 255270
rect 352564 255206 352616 255212
rect 300124 203788 300176 203794
rect 300124 203730 300176 203736
rect 364996 203658 365024 425206
rect 429212 424386 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 427378 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 497554 477540 702406
rect 477500 497548 477552 497554
rect 477500 497490 477552 497496
rect 462320 427372 462372 427378
rect 462320 427314 462372 427320
rect 494072 424658 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 453354 527220 703520
rect 543476 700534 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 535736 700528 535788 700534
rect 535736 700470 535788 700476
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 534356 696992 534408 696998
rect 534356 696934 534408 696940
rect 534172 630692 534224 630698
rect 534172 630634 534224 630640
rect 533344 616888 533396 616894
rect 533344 616830 533396 616836
rect 532884 590708 532936 590714
rect 532884 590650 532936 590656
rect 532792 576904 532844 576910
rect 532792 576846 532844 576852
rect 531320 524476 531372 524482
rect 531320 524418 531372 524424
rect 530124 484424 530176 484430
rect 530124 484366 530176 484372
rect 527180 453348 527232 453354
rect 527180 453290 527232 453296
rect 529664 430636 529716 430642
rect 529664 430578 529716 430584
rect 494060 424652 494112 424658
rect 494060 424594 494112 424600
rect 445024 424448 445076 424454
rect 445024 424390 445076 424396
rect 429200 424380 429252 424386
rect 429200 424322 429252 424328
rect 429212 420102 429240 424322
rect 444930 420336 444986 420345
rect 444930 420271 444986 420280
rect 444746 420200 444802 420209
rect 444746 420135 444802 420144
rect 429200 420096 429252 420102
rect 429200 420038 429252 420044
rect 444760 346390 444788 420135
rect 444748 346384 444800 346390
rect 444748 346326 444800 346332
rect 444944 293962 444972 420271
rect 444932 293956 444984 293962
rect 444932 293898 444984 293904
rect 440884 244928 440936 244934
rect 440884 244870 440936 244876
rect 440896 224262 440924 244870
rect 440884 224256 440936 224262
rect 440884 224198 440936 224204
rect 364984 203652 365036 203658
rect 364984 203594 365036 203600
rect 284944 202564 284996 202570
rect 284944 202506 284996 202512
rect 445036 202502 445064 424390
rect 529204 424380 529256 424386
rect 529204 424322 529256 424328
rect 445300 423292 445352 423298
rect 445300 423234 445352 423240
rect 445116 423224 445168 423230
rect 445116 423166 445168 423172
rect 445024 202496 445076 202502
rect 445024 202438 445076 202444
rect 445128 202434 445156 423166
rect 445208 422680 445260 422686
rect 445208 422622 445260 422628
rect 445116 202428 445168 202434
rect 445116 202370 445168 202376
rect 445220 202366 445248 422622
rect 445208 202360 445260 202366
rect 445208 202302 445260 202308
rect 445312 202298 445340 423234
rect 524144 423156 524196 423162
rect 524144 423098 524196 423104
rect 445390 422920 445446 422929
rect 445390 422855 445446 422864
rect 522948 422884 523000 422890
rect 445404 202842 445432 422855
rect 522948 422826 523000 422832
rect 522028 422816 522080 422822
rect 522028 422758 522080 422764
rect 521016 421320 521068 421326
rect 521016 421262 521068 421268
rect 520648 421184 520700 421190
rect 520648 421126 520700 421132
rect 445574 420064 445630 420073
rect 445574 419999 445630 420008
rect 445484 419892 445536 419898
rect 445484 419834 445536 419840
rect 445392 202836 445444 202842
rect 445392 202778 445444 202784
rect 445300 202292 445352 202298
rect 445300 202234 445352 202240
rect 256056 202224 256108 202230
rect 256056 202166 256108 202172
rect 256068 201550 256096 202166
rect 261576 201680 261628 201686
rect 261576 201622 261628 201628
rect 260104 201612 260156 201618
rect 260104 201554 260156 201560
rect 256056 201544 256108 201550
rect 256056 201486 256108 201492
rect 251364 200932 251416 200938
rect 251364 200874 251416 200880
rect 246580 200864 246632 200870
rect 246580 200806 246632 200812
rect 241888 200796 241940 200802
rect 241888 200738 241940 200744
rect 241900 200462 241928 200738
rect 241888 200456 241940 200462
rect 241888 200398 241940 200404
rect 241900 199866 241928 200398
rect 246592 200394 246620 200806
rect 246580 200388 246632 200394
rect 246580 200330 246632 200336
rect 246592 199866 246620 200330
rect 251376 200326 251404 200874
rect 251364 200320 251416 200326
rect 251364 200262 251416 200268
rect 251376 199866 251404 200262
rect 256068 199866 256096 201486
rect 222488 199838 222916 199866
rect 227180 199838 227608 199866
rect 231964 199838 232392 199866
rect 236656 199838 237084 199866
rect 241868 199838 241928 199866
rect 246560 199838 246620 199866
rect 251344 199838 251404 199866
rect 256036 199838 256096 199866
rect 185012 199702 185072 199730
rect 218132 199702 218192 199730
rect 79324 137964 79376 137970
rect 79324 137906 79376 137912
rect 260116 126954 260144 201554
rect 261484 200524 261536 200530
rect 261484 200466 261536 200472
rect 260104 126948 260156 126954
rect 260104 126890 260156 126896
rect 77944 85536 77996 85542
rect 77944 85478 77996 85484
rect 80118 79914 80146 80036
rect 79980 79886 80146 79914
rect 79980 79694 80008 79886
rect 80060 79824 80112 79830
rect 80060 79766 80112 79772
rect 80152 79824 80204 79830
rect 80152 79766 80204 79772
rect 79968 79688 80020 79694
rect 79968 79630 80020 79636
rect 70400 78532 70452 78538
rect 70400 78474 70452 78480
rect 65524 78464 65576 78470
rect 65524 78406 65576 78412
rect 53104 78396 53156 78402
rect 53104 78338 53156 78344
rect 50344 78328 50396 78334
rect 50344 78270 50396 78276
rect 28264 78260 28316 78266
rect 28264 78202 28316 78208
rect 25504 78124 25556 78130
rect 25504 78066 25556 78072
rect 15844 78056 15896 78062
rect 15844 77998 15896 78004
rect 10324 77988 10376 77994
rect 10324 77930 10376 77936
rect 3790 32464 3846 32473
rect 3790 32399 3846 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 3608 10328 3660 10334
rect 3608 10270 3660 10276
rect 2872 7608 2924 7614
rect 2872 7550 2924 7556
rect 2884 480 2912 7550
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 542 -960 654 326
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 3620 354 3648 10270
rect 7656 7676 7708 7682
rect 7656 7618 7708 7624
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5276 480 5304 3470
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 7618
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8772 480 8800 6122
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 14418
rect 10336 3534 10364 77930
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15212 16574 15240 17206
rect 15212 16546 15792 16574
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 13544 10396 13596 10402
rect 13544 10338 13596 10344
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 11164 480 11192 3538
rect 12360 480 12388 4762
rect 13556 480 13584 10338
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 14486
rect 15764 3482 15792 16546
rect 15856 3602 15884 77998
rect 22100 43444 22152 43450
rect 22100 43386 22152 43392
rect 16580 42152 16632 42158
rect 16580 42094 16632 42100
rect 16592 16574 16620 42094
rect 22112 16574 22140 43386
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24872 16574 24900 18566
rect 16592 16546 17080 16574
rect 22112 16546 22600 16574
rect 24872 16546 25360 16574
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15764 3454 15976 3482
rect 15948 480 15976 3454
rect 17052 480 17080 16546
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 11698
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 480 19472 2994
rect 20640 480 20668 3606
rect 21836 480 21864 7686
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24216 15904 24268 15910
rect 24216 15846 24268 15852
rect 24228 480 24256 15846
rect 25332 480 25360 16546
rect 25516 3058 25544 78066
rect 27712 13116 27764 13122
rect 27712 13058 27764 13064
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 26528 480 26556 8910
rect 27724 480 27752 13058
rect 28276 3670 28304 78202
rect 32404 78192 32456 78198
rect 32404 78134 32456 78140
rect 30380 44872 30432 44878
rect 30380 44814 30432 44820
rect 30392 16574 30420 44814
rect 30392 16546 30880 16574
rect 30104 9036 30156 9042
rect 30104 8978 30156 8984
rect 28264 3664 28316 3670
rect 28264 3606 28316 3612
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 28920 480 28948 3470
rect 30116 480 30144 8978
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31944 15972 31996 15978
rect 31944 15914 31996 15920
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 15914
rect 32416 3534 32444 78134
rect 49700 76560 49752 76566
rect 49700 76502 49752 76508
rect 37280 75200 37332 75206
rect 37280 75142 37332 75148
rect 35900 42220 35952 42226
rect 35900 42162 35952 42168
rect 35912 16574 35940 42162
rect 37292 16574 37320 75142
rect 44180 40792 44232 40798
rect 44180 40734 44232 40740
rect 38660 17332 38712 17338
rect 38660 17274 38712 17280
rect 38672 16574 38700 17274
rect 35912 16546 36768 16574
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 34520 13184 34572 13190
rect 34520 13126 34572 13132
rect 33600 6248 33652 6254
rect 33600 6190 33652 6196
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33612 480 33640 6190
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 13126
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 36004 480 36032 3334
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 41880 13252 41932 13258
rect 41880 13194 41932 13200
rect 40224 10464 40276 10470
rect 40224 10406 40276 10412
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 10406
rect 41892 480 41920 13194
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 43088 480 43116 3538
rect 44192 3534 44220 40734
rect 45560 17400 45612 17406
rect 45560 17342 45612 17348
rect 45572 16574 45600 17342
rect 49712 16574 49740 76502
rect 45572 16546 46704 16574
rect 49712 16546 50200 16574
rect 44272 11824 44324 11830
rect 44272 11766 44324 11772
rect 44180 3528 44232 3534
rect 44180 3470 44232 3476
rect 44284 480 44312 11766
rect 45100 3528 45152 3534
rect 45100 3470 45152 3476
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45112 354 45140 3470
rect 46676 480 46704 16546
rect 47860 7812 47912 7818
rect 47860 7754 47912 7760
rect 47872 480 47900 7754
rect 48964 6316 49016 6322
rect 48964 6258 49016 6264
rect 48976 480 49004 6258
rect 50172 480 50200 16546
rect 50356 3534 50384 78270
rect 51080 76628 51132 76634
rect 51080 76570 51132 76576
rect 50344 3528 50396 3534
rect 50344 3470 50396 3476
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 76570
rect 52460 49020 52512 49026
rect 52460 48962 52512 48968
rect 52472 16574 52500 48962
rect 52472 16546 52592 16574
rect 52564 480 52592 16546
rect 53012 14612 53064 14618
rect 53012 14554 53064 14560
rect 53024 490 53052 14554
rect 53116 3602 53144 78338
rect 59360 43512 59412 43518
rect 59360 43454 59412 43460
rect 53840 22772 53892 22778
rect 53840 22714 53892 22720
rect 53852 16574 53880 22714
rect 53852 16546 54984 16574
rect 53104 3596 53156 3602
rect 53104 3538 53156 3544
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53024 462 53328 490
rect 54956 480 54984 16546
rect 56784 14680 56836 14686
rect 56784 14622 56836 14628
rect 56048 10532 56100 10538
rect 56048 10474 56100 10480
rect 56060 480 56088 10474
rect 53300 354 53328 462
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 14622
rect 58440 9104 58492 9110
rect 58440 9046 58492 9052
rect 58452 480 58480 9046
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 43454
rect 60740 17468 60792 17474
rect 60740 17410 60792 17416
rect 60752 16574 60780 17410
rect 60752 16546 60872 16574
rect 60844 480 60872 16546
rect 61568 11960 61620 11966
rect 61568 11902 61620 11908
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 11902
rect 63224 11892 63276 11898
rect 63224 11834 63276 11840
rect 63236 480 63264 11834
rect 65536 4146 65564 78406
rect 66260 43580 66312 43586
rect 66260 43522 66312 43528
rect 66272 16574 66300 43522
rect 70412 16574 70440 78474
rect 73160 43648 73212 43654
rect 73160 43590 73212 43596
rect 73172 16574 73200 43590
rect 77300 21412 77352 21418
rect 77300 21354 77352 21360
rect 77312 16574 77340 21354
rect 66272 16546 66760 16574
rect 70412 16546 71544 16574
rect 73172 16546 73384 16574
rect 77312 16546 78168 16574
rect 65616 4888 65668 4894
rect 65616 4830 65668 4836
rect 64328 4140 64380 4146
rect 64328 4082 64380 4088
rect 65524 4140 65576 4146
rect 65524 4082 65576 4088
rect 64340 480 64368 4082
rect 65628 2530 65656 4830
rect 65536 2502 65656 2530
rect 65536 480 65564 2502
rect 66732 480 66760 16546
rect 67640 16040 67692 16046
rect 67640 15982 67692 15988
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 15982
rect 69848 13320 69900 13326
rect 69848 13262 69900 13268
rect 69112 4956 69164 4962
rect 69112 4898 69164 4904
rect 69124 480 69152 4898
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 13262
rect 71516 480 71544 16546
rect 72608 9172 72660 9178
rect 72608 9114 72660 9120
rect 72620 480 72648 9114
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75000 16108 75052 16114
rect 75000 16050 75052 16056
rect 75012 480 75040 16050
rect 77392 6384 77444 6390
rect 77392 6326 77444 6332
rect 76196 5024 76248 5030
rect 76196 4966 76248 4972
rect 76208 480 76236 4966
rect 77404 480 77432 6326
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 80072 7614 80100 79766
rect 80164 10334 80192 79766
rect 80244 79688 80296 79694
rect 80394 79642 80422 80036
rect 80762 79898 80790 80036
rect 80750 79892 80802 79898
rect 80750 79834 80802 79840
rect 81130 79830 81158 80036
rect 81498 79914 81526 80036
rect 81452 79886 81526 79914
rect 81118 79824 81170 79830
rect 81118 79766 81170 79772
rect 80244 79630 80296 79636
rect 80256 78742 80284 79630
rect 80348 79614 80422 79642
rect 80348 78810 80376 79614
rect 80336 78804 80388 78810
rect 80336 78746 80388 78752
rect 80244 78736 80296 78742
rect 80244 78678 80296 78684
rect 80256 40730 80284 78678
rect 80348 42090 80376 78746
rect 81452 77994 81480 79886
rect 81624 79824 81676 79830
rect 81866 79778 81894 80036
rect 82234 79830 82262 80036
rect 81624 79766 81676 79772
rect 81440 77988 81492 77994
rect 81440 77930 81492 77936
rect 81532 77308 81584 77314
rect 81532 77250 81584 77256
rect 80336 42084 80388 42090
rect 80336 42026 80388 42032
rect 80244 40724 80296 40730
rect 80244 40666 80296 40672
rect 80152 10328 80204 10334
rect 80152 10270 80204 10276
rect 80060 7608 80112 7614
rect 80060 7550 80112 7556
rect 80888 7608 80940 7614
rect 80888 7550 80940 7556
rect 79692 5092 79744 5098
rect 79692 5034 79744 5040
rect 79704 480 79732 5034
rect 80900 480 80928 7550
rect 81544 6186 81572 77250
rect 81636 7682 81664 79766
rect 81820 79750 81894 79778
rect 82222 79824 82274 79830
rect 82602 79778 82630 80036
rect 82222 79766 82274 79772
rect 82556 79750 82630 79778
rect 82976 79778 83004 80036
rect 83338 79914 83366 80036
rect 83292 79886 83366 79914
rect 82976 79750 83044 79778
rect 81624 7676 81676 7682
rect 81624 7618 81676 7624
rect 81532 6180 81584 6186
rect 81532 6122 81584 6128
rect 81820 3466 81848 79750
rect 82556 77314 82584 79750
rect 82544 77308 82596 77314
rect 82544 77250 82596 77256
rect 82912 77308 82964 77314
rect 82912 77250 82964 77256
rect 82924 10402 82952 77250
rect 83016 14482 83044 79750
rect 83292 78062 83320 79886
rect 83706 79778 83734 80036
rect 84074 79778 84102 80036
rect 84442 79778 84470 80036
rect 84810 79778 84838 80036
rect 85178 79778 85206 80036
rect 83476 79750 83734 79778
rect 84028 79750 84102 79778
rect 84212 79750 84470 79778
rect 84580 79750 84838 79778
rect 84948 79750 85206 79778
rect 85552 79778 85580 80036
rect 85920 79778 85948 80036
rect 86282 79778 86310 80036
rect 86650 79778 86678 80036
rect 87018 79778 87046 80036
rect 87386 79778 87414 80036
rect 87754 79778 87782 80036
rect 88122 79778 88150 80036
rect 88490 79778 88518 80036
rect 88858 79914 88886 80036
rect 85552 79750 85712 79778
rect 85920 79750 85988 79778
rect 83280 78056 83332 78062
rect 83280 77998 83332 78004
rect 83476 64874 83504 79750
rect 84028 77314 84056 79750
rect 84016 77308 84068 77314
rect 84016 77250 84068 77256
rect 83108 64846 83504 64874
rect 83004 14476 83056 14482
rect 83004 14418 83056 14424
rect 82912 10396 82964 10402
rect 82912 10338 82964 10344
rect 82084 7880 82136 7886
rect 82084 7822 82136 7828
rect 81808 3460 81860 3466
rect 81808 3402 81860 3408
rect 82096 480 82124 7822
rect 83108 4826 83136 64846
rect 84212 14550 84240 79750
rect 84580 77296 84608 79750
rect 84304 77268 84608 77296
rect 84304 17270 84332 77268
rect 84948 64874 84976 79750
rect 84396 64846 84976 64874
rect 84396 42158 84424 64846
rect 84384 42152 84436 42158
rect 84384 42094 84436 42100
rect 84292 17264 84344 17270
rect 84292 17206 84344 17212
rect 84200 14544 84252 14550
rect 84200 14486 84252 14492
rect 85684 11762 85712 79750
rect 85960 78130 85988 79750
rect 86236 79750 86310 79778
rect 86420 79750 86678 79778
rect 86972 79750 87046 79778
rect 87156 79750 87414 79778
rect 87708 79750 87782 79778
rect 88076 79750 88150 79778
rect 88444 79750 88518 79778
rect 88812 79886 88886 79914
rect 86236 78266 86264 79750
rect 86224 78260 86276 78266
rect 86224 78202 86276 78208
rect 85948 78124 86000 78130
rect 85948 78066 86000 78072
rect 86420 64874 86448 79750
rect 86972 77314 87000 79750
rect 86960 77308 87012 77314
rect 87156 77296 87184 79750
rect 86960 77250 87012 77256
rect 87064 77268 87184 77296
rect 87236 77308 87288 77314
rect 86960 75676 87012 75682
rect 86960 75618 87012 75624
rect 85868 64846 86448 64874
rect 85764 14476 85816 14482
rect 85764 14418 85816 14424
rect 85672 11756 85724 11762
rect 85672 11698 85724 11704
rect 85776 6914 85804 14418
rect 85868 7750 85896 64846
rect 86868 9240 86920 9246
rect 86868 9182 86920 9188
rect 85856 7744 85908 7750
rect 85856 7686 85908 7692
rect 85684 6886 85804 6914
rect 84476 6180 84528 6186
rect 84476 6122 84528 6128
rect 83280 5160 83332 5166
rect 83280 5102 83332 5108
rect 83096 4820 83148 4826
rect 83096 4762 83148 4768
rect 83292 480 83320 5102
rect 84488 480 84516 6122
rect 85684 480 85712 6886
rect 86880 480 86908 9182
rect 86972 8974 87000 75618
rect 87064 15910 87092 77268
rect 87236 77250 87288 77256
rect 87144 77172 87196 77178
rect 87144 77114 87196 77120
rect 87156 18630 87184 77114
rect 87248 43450 87276 77250
rect 87708 77178 87736 79750
rect 87696 77172 87748 77178
rect 87696 77114 87748 77120
rect 88076 75682 88104 79750
rect 88064 75676 88116 75682
rect 88064 75618 88116 75624
rect 87236 43444 87288 43450
rect 87236 43386 87288 43392
rect 87144 18624 87196 18630
rect 87144 18566 87196 18572
rect 87052 15904 87104 15910
rect 87052 15846 87104 15852
rect 88444 13122 88472 79750
rect 88812 78198 88840 79886
rect 89226 79778 89254 80036
rect 89594 79778 89622 80036
rect 89812 79892 89864 79898
rect 89812 79834 89864 79840
rect 88996 79750 89254 79778
rect 89548 79750 89622 79778
rect 89720 79824 89772 79830
rect 89720 79766 89772 79772
rect 88800 78192 88852 78198
rect 88800 78134 88852 78140
rect 88524 77308 88576 77314
rect 88524 77250 88576 77256
rect 88536 44878 88564 77250
rect 88996 64874 89024 79750
rect 89548 77314 89576 79750
rect 89536 77308 89588 77314
rect 89536 77250 89588 77256
rect 88628 64846 89024 64874
rect 88524 44872 88576 44878
rect 88524 44814 88576 44820
rect 88432 13116 88484 13122
rect 88432 13058 88484 13064
rect 87512 10328 87564 10334
rect 87512 10270 87564 10276
rect 86960 8968 87012 8974
rect 86960 8910 87012 8916
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 10270
rect 88628 9042 88656 64846
rect 89168 11756 89220 11762
rect 89168 11698 89220 11704
rect 88616 9036 88668 9042
rect 88616 8978 88668 8984
rect 89180 480 89208 11698
rect 89732 6254 89760 79766
rect 89824 13190 89852 79834
rect 89962 79778 89990 80036
rect 90330 79830 90358 80036
rect 90698 79898 90726 80036
rect 90686 79892 90738 79898
rect 90686 79834 90738 79840
rect 89916 79750 89990 79778
rect 90318 79824 90370 79830
rect 90318 79766 90370 79772
rect 91072 79778 91100 80036
rect 91434 79778 91462 80036
rect 91802 79914 91830 80036
rect 91072 79750 91140 79778
rect 89916 15978 89944 79750
rect 91112 78334 91140 79750
rect 91204 79750 91462 79778
rect 91756 79886 91830 79914
rect 91100 78328 91152 78334
rect 91100 78270 91152 78276
rect 91204 42226 91232 79750
rect 91756 75206 91784 79886
rect 92078 79778 92106 80036
rect 91848 79750 92106 79778
rect 92452 79778 92480 80036
rect 92820 79778 92848 80036
rect 93188 79778 93216 80036
rect 93550 79778 93578 80036
rect 92452 79750 92704 79778
rect 92820 79750 92888 79778
rect 93188 79750 93256 79778
rect 91744 75200 91796 75206
rect 91744 75142 91796 75148
rect 91848 60734 91876 79750
rect 92676 77602 92704 79750
rect 92676 77574 92796 77602
rect 92572 77172 92624 77178
rect 92572 77114 92624 77120
rect 91296 60706 91876 60734
rect 91192 42220 91244 42226
rect 91192 42162 91244 42168
rect 91296 17338 91324 60706
rect 91284 17332 91336 17338
rect 91284 17274 91336 17280
rect 89904 15972 89956 15978
rect 89904 15914 89956 15920
rect 89812 13184 89864 13190
rect 89812 13126 89864 13132
rect 92584 11830 92612 77114
rect 92768 65618 92796 77574
rect 92756 65612 92808 65618
rect 92756 65554 92808 65560
rect 92756 65408 92808 65414
rect 92756 65350 92808 65356
rect 92664 58608 92716 58614
rect 92664 58550 92716 58556
rect 92676 13258 92704 58550
rect 92664 13252 92716 13258
rect 92664 13194 92716 13200
rect 92572 11824 92624 11830
rect 92572 11766 92624 11772
rect 92768 10470 92796 65350
rect 92860 58614 92888 79750
rect 93228 78402 93256 79750
rect 93504 79750 93578 79778
rect 93924 79778 93952 80036
rect 94286 79778 94314 80036
rect 94654 79778 94682 80036
rect 95022 79778 95050 80036
rect 95390 79914 95418 80036
rect 95758 79914 95786 80036
rect 93924 79750 93992 79778
rect 93216 78396 93268 78402
rect 93216 78338 93268 78344
rect 93124 78328 93176 78334
rect 93124 78270 93176 78276
rect 92848 58608 92900 58614
rect 92848 58550 92900 58556
rect 93136 14618 93164 78270
rect 93504 77178 93532 79750
rect 93964 77314 93992 79750
rect 94056 79750 94314 79778
rect 94608 79750 94682 79778
rect 94976 79750 95050 79778
rect 95344 79886 95418 79914
rect 95712 79886 95786 79914
rect 93952 77308 94004 77314
rect 93952 77250 94004 77256
rect 93860 77240 93912 77246
rect 93860 77182 93912 77188
rect 93492 77172 93544 77178
rect 93492 77114 93544 77120
rect 93124 14612 93176 14618
rect 93124 14554 93176 14560
rect 92756 10464 92808 10470
rect 92756 10406 92808 10412
rect 92572 10396 92624 10402
rect 92572 10338 92624 10344
rect 90364 7676 90416 7682
rect 90364 7618 90416 7624
rect 89720 6248 89772 6254
rect 89720 6190 89772 6196
rect 90376 480 90404 7618
rect 91560 6248 91612 6254
rect 91560 6190 91612 6196
rect 91572 480 91600 6190
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92584 354 92612 10338
rect 93872 6322 93900 77182
rect 93952 77172 94004 77178
rect 93952 77114 94004 77120
rect 93964 7818 93992 77114
rect 94056 17406 94084 79750
rect 94136 77308 94188 77314
rect 94136 77250 94188 77256
rect 94148 40798 94176 77250
rect 94608 77178 94636 79750
rect 94976 77246 95004 79750
rect 94964 77240 95016 77246
rect 94964 77182 95016 77188
rect 94596 77172 94648 77178
rect 94596 77114 94648 77120
rect 95344 76566 95372 79886
rect 95712 76634 95740 79886
rect 96126 79778 96154 80036
rect 96494 79778 96522 80036
rect 96712 79892 96764 79898
rect 96712 79834 96764 79840
rect 95988 79750 96154 79778
rect 96448 79750 96522 79778
rect 96620 79824 96672 79830
rect 96620 79766 96672 79772
rect 95700 76628 95752 76634
rect 95700 76570 95752 76576
rect 95332 76560 95384 76566
rect 95332 76502 95384 76508
rect 95988 60734 96016 79750
rect 96448 78334 96476 79750
rect 96436 78328 96488 78334
rect 96436 78270 96488 78276
rect 95436 60706 96016 60734
rect 95436 49026 95464 60706
rect 95424 49020 95476 49026
rect 95424 48962 95476 48968
rect 94228 40928 94280 40934
rect 94228 40870 94280 40876
rect 94136 40792 94188 40798
rect 94136 40734 94188 40740
rect 94044 17400 94096 17406
rect 94044 17342 94096 17348
rect 94240 16574 94268 40870
rect 94240 16546 94728 16574
rect 93952 7812 94004 7818
rect 93952 7754 94004 7760
rect 93860 6316 93912 6322
rect 93860 6258 93912 6264
rect 93952 3392 94004 3398
rect 93952 3334 94004 3340
rect 93964 480 93992 3334
rect 92726 354 92838 480
rect 92584 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 96632 10538 96660 79766
rect 96724 14686 96752 79834
rect 96862 79778 96890 80036
rect 97230 79830 97258 80036
rect 97598 79898 97626 80036
rect 97586 79892 97638 79898
rect 97586 79834 97638 79840
rect 96816 79750 96890 79778
rect 97218 79824 97270 79830
rect 97218 79766 97270 79772
rect 97972 79778 98000 80036
rect 98092 79892 98144 79898
rect 98092 79834 98144 79840
rect 97972 79750 98040 79778
rect 96816 22778 96844 79750
rect 97264 78600 97316 78606
rect 97264 78542 97316 78548
rect 96804 22772 96856 22778
rect 96804 22714 96856 22720
rect 96712 14680 96764 14686
rect 96712 14622 96764 14628
rect 96620 10532 96672 10538
rect 96620 10474 96672 10480
rect 97276 7886 97304 78542
rect 98012 9110 98040 79750
rect 98104 11966 98132 79834
rect 98184 79824 98236 79830
rect 98334 79778 98362 80036
rect 98702 79830 98730 80036
rect 99070 79898 99098 80036
rect 99058 79892 99110 79898
rect 99058 79834 99110 79840
rect 98184 79766 98236 79772
rect 98196 17474 98224 79766
rect 98288 79750 98362 79778
rect 98690 79824 98742 79830
rect 98690 79766 98742 79772
rect 99444 79778 99472 80036
rect 99806 79914 99834 80036
rect 99760 79886 99834 79914
rect 99564 79824 99616 79830
rect 99444 79750 99512 79778
rect 99564 79766 99616 79772
rect 98288 43518 98316 79750
rect 98276 43512 98328 43518
rect 98276 43454 98328 43460
rect 98276 19984 98328 19990
rect 98276 19926 98328 19932
rect 98184 17468 98236 17474
rect 98184 17410 98236 17416
rect 98092 11960 98144 11966
rect 98092 11902 98144 11908
rect 98000 9104 98052 9110
rect 98000 9046 98052 9052
rect 97264 7880 97316 7886
rect 97264 7822 97316 7828
rect 97448 7744 97500 7750
rect 97448 7686 97500 7692
rect 96252 3324 96304 3330
rect 96252 3266 96304 3272
rect 96264 480 96292 3266
rect 97460 480 97488 7686
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98288 354 98316 19926
rect 99484 11898 99512 79750
rect 99576 43586 99604 79766
rect 99760 78470 99788 79886
rect 100174 79778 100202 80036
rect 100542 79830 100570 80036
rect 99944 79750 100202 79778
rect 100530 79824 100582 79830
rect 100530 79766 100582 79772
rect 100916 79778 100944 80036
rect 101278 79778 101306 80036
rect 101646 79778 101674 80036
rect 102014 79778 102042 80036
rect 102382 79778 102410 80036
rect 102750 79778 102778 80036
rect 103118 79778 103146 80036
rect 100916 79750 100984 79778
rect 99748 78464 99800 78470
rect 99748 78406 99800 78412
rect 99944 64874 99972 79750
rect 100024 77376 100076 77382
rect 100024 77318 100076 77324
rect 99668 64846 99972 64874
rect 99564 43580 99616 43586
rect 99564 43522 99616 43528
rect 99472 11892 99524 11898
rect 99472 11834 99524 11840
rect 99668 4894 99696 64846
rect 100036 16114 100064 77318
rect 100852 77308 100904 77314
rect 100852 77250 100904 77256
rect 100024 16108 100076 16114
rect 100024 16050 100076 16056
rect 100864 13326 100892 77250
rect 100956 16046 100984 79750
rect 101048 79750 101306 79778
rect 101600 79750 101674 79778
rect 101968 79750 102042 79778
rect 102244 79750 102410 79778
rect 102612 79750 102778 79778
rect 103072 79750 103146 79778
rect 103492 79778 103520 80036
rect 103612 79824 103664 79830
rect 103492 79750 103560 79778
rect 103854 79778 103882 80036
rect 104130 79778 104158 80036
rect 104498 79830 104526 80036
rect 103612 79766 103664 79772
rect 100944 16040 100996 16046
rect 100944 15982 100996 15988
rect 100852 13320 100904 13326
rect 100852 13262 100904 13268
rect 101048 11778 101076 79750
rect 101404 78124 101456 78130
rect 101404 78066 101456 78072
rect 101416 14482 101444 78066
rect 101600 77314 101628 79750
rect 101968 78538 101996 79750
rect 101956 78532 102008 78538
rect 101956 78474 102008 78480
rect 102140 77988 102192 77994
rect 102140 77930 102192 77936
rect 101588 77308 101640 77314
rect 101588 77250 101640 77256
rect 101404 14476 101456 14482
rect 101404 14418 101456 14424
rect 100956 11750 101076 11778
rect 100956 4962 100984 11750
rect 101036 8968 101088 8974
rect 101036 8910 101088 8916
rect 100944 4956 100996 4962
rect 100944 4898 100996 4904
rect 99656 4888 99708 4894
rect 99656 4830 99708 4836
rect 99840 3596 99892 3602
rect 99840 3538 99892 3544
rect 99852 480 99880 3538
rect 101048 480 101076 8910
rect 102152 3534 102180 77930
rect 102244 9178 102272 79750
rect 102612 64874 102640 79750
rect 103072 77382 103100 79750
rect 103060 77376 103112 77382
rect 103060 77318 103112 77324
rect 102336 64846 102640 64874
rect 102336 43654 102364 64846
rect 102324 43648 102376 43654
rect 102324 43590 102376 43596
rect 102324 43444 102376 43450
rect 102324 43386 102376 43392
rect 102232 9172 102284 9178
rect 102232 9114 102284 9120
rect 102336 6914 102364 43386
rect 102244 6886 102364 6914
rect 102140 3528 102192 3534
rect 102140 3470 102192 3476
rect 102244 480 102272 6886
rect 103532 5030 103560 79750
rect 103624 5098 103652 79766
rect 103716 79750 103882 79778
rect 103992 79750 104158 79778
rect 104486 79824 104538 79830
rect 104486 79766 104538 79772
rect 104872 79778 104900 80036
rect 105240 79914 105268 80036
rect 105240 79886 105308 79914
rect 104872 79750 105124 79778
rect 103716 6390 103744 79750
rect 103992 64874 104020 79750
rect 104992 77308 105044 77314
rect 104992 77250 105044 77256
rect 103808 64846 104020 64874
rect 103808 21418 103836 64846
rect 103888 22160 103940 22166
rect 103888 22102 103940 22108
rect 103796 21412 103848 21418
rect 103796 21354 103848 21360
rect 103900 16574 103928 22102
rect 103900 16546 104112 16574
rect 103704 6384 103756 6390
rect 103704 6326 103756 6332
rect 103612 5092 103664 5098
rect 103612 5034 103664 5040
rect 103520 5024 103572 5030
rect 103520 4966 103572 4972
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 103428 3528 103480 3534
rect 103428 3470 103480 3476
rect 103348 480 103376 3470
rect 103440 3330 103468 3470
rect 103428 3324 103480 3330
rect 103428 3266 103480 3272
rect 98614 354 98726 480
rect 98288 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105004 6186 105032 77250
rect 105096 7614 105124 79750
rect 105280 78606 105308 79886
rect 105602 79778 105630 80036
rect 105970 79778 105998 80036
rect 106338 79914 106366 80036
rect 105464 79750 105630 79778
rect 105924 79750 105998 79778
rect 106292 79886 106366 79914
rect 105268 78600 105320 78606
rect 105268 78542 105320 78548
rect 105464 64874 105492 79750
rect 105544 77444 105596 77450
rect 105544 77386 105596 77392
rect 105188 64846 105492 64874
rect 105084 7608 105136 7614
rect 105084 7550 105136 7556
rect 104992 6180 105044 6186
rect 104992 6122 105044 6128
rect 105188 5166 105216 64846
rect 105556 11762 105584 77386
rect 105924 77314 105952 79750
rect 106292 78130 106320 79886
rect 106372 79824 106424 79830
rect 106706 79778 106734 80036
rect 107074 79830 107102 80036
rect 106372 79766 106424 79772
rect 106280 78124 106332 78130
rect 106280 78066 106332 78072
rect 105912 77308 105964 77314
rect 105912 77250 105964 77256
rect 105544 11756 105596 11762
rect 105544 11698 105596 11704
rect 106384 10334 106412 79766
rect 106476 79750 106734 79778
rect 107062 79824 107114 79830
rect 107442 79778 107470 80036
rect 107062 79766 107114 79772
rect 107396 79750 107470 79778
rect 107816 79778 107844 80036
rect 108178 79778 108206 80036
rect 108546 79778 108574 80036
rect 108914 79778 108942 80036
rect 109282 79778 109310 80036
rect 109650 79914 109678 80036
rect 107816 79750 107884 79778
rect 106372 10328 106424 10334
rect 106372 10270 106424 10276
rect 106476 9246 106504 79750
rect 106924 77512 106976 77518
rect 106924 77454 106976 77460
rect 106464 9240 106516 9246
rect 106464 9182 106516 9188
rect 106936 6914 106964 77454
rect 107396 77450 107424 79750
rect 107660 77852 107712 77858
rect 107660 77794 107712 77800
rect 107384 77444 107436 77450
rect 107384 77386 107436 77392
rect 107016 77376 107068 77382
rect 107016 77318 107068 77324
rect 107028 10402 107056 77318
rect 107016 10396 107068 10402
rect 107016 10338 107068 10344
rect 106844 6886 106964 6914
rect 105176 5160 105228 5166
rect 105176 5102 105228 5108
rect 105728 4208 105780 4214
rect 105728 4150 105780 4156
rect 105740 480 105768 4150
rect 106844 3466 106872 6886
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107672 3482 107700 77794
rect 107752 77308 107804 77314
rect 107752 77250 107804 77256
rect 107764 6254 107792 77250
rect 107856 7682 107884 79750
rect 108132 79750 108206 79778
rect 108500 79750 108574 79778
rect 108868 79750 108942 79778
rect 109144 79750 109310 79778
rect 109604 79886 109678 79914
rect 108132 77314 108160 79750
rect 108500 77382 108528 79750
rect 108868 77518 108896 79750
rect 108856 77512 108908 77518
rect 108856 77454 108908 77460
rect 108488 77376 108540 77382
rect 108488 77318 108540 77324
rect 108120 77308 108172 77314
rect 108120 77250 108172 77256
rect 108304 77308 108356 77314
rect 108304 77250 108356 77256
rect 107844 7676 107896 7682
rect 107844 7618 107896 7624
rect 107752 6248 107804 6254
rect 107752 6190 107804 6196
rect 108316 3602 108344 77250
rect 109144 40934 109172 79750
rect 109604 77314 109632 79886
rect 110018 79778 110046 80036
rect 109972 79750 110046 79778
rect 110392 79778 110420 80036
rect 110754 79914 110782 80036
rect 111122 79914 111150 80036
rect 110708 79886 110782 79914
rect 111076 79886 111150 79914
rect 110392 79750 110644 79778
rect 109592 77308 109644 77314
rect 109592 77250 109644 77256
rect 109684 77308 109736 77314
rect 109684 77250 109736 77256
rect 109224 77240 109276 77246
rect 109224 77182 109276 77188
rect 109132 40928 109184 40934
rect 109132 40870 109184 40876
rect 109236 7750 109264 77182
rect 109224 7744 109276 7750
rect 109224 7686 109276 7692
rect 109696 3670 109724 77250
rect 109972 77246 110000 79750
rect 110420 78396 110472 78402
rect 110420 78338 110472 78344
rect 109960 77240 110012 77246
rect 109960 77182 110012 77188
rect 110432 6914 110460 78338
rect 110512 78260 110564 78266
rect 110512 78202 110564 78208
rect 110524 8974 110552 78202
rect 110616 19990 110644 79750
rect 110708 77314 110736 79886
rect 111076 78266 111104 79886
rect 111490 79778 111518 80036
rect 111858 79914 111886 80036
rect 111444 79750 111518 79778
rect 111812 79886 111886 79914
rect 111064 78260 111116 78266
rect 111064 78202 111116 78208
rect 111064 78124 111116 78130
rect 111064 78066 111116 78072
rect 110696 77308 110748 77314
rect 110696 77250 110748 77256
rect 110696 77172 110748 77178
rect 110696 77114 110748 77120
rect 110708 43450 110736 77114
rect 110696 43444 110748 43450
rect 110696 43386 110748 43392
rect 110696 23452 110748 23458
rect 110696 23394 110748 23400
rect 110604 19984 110656 19990
rect 110604 19926 110656 19932
rect 110708 16574 110736 23394
rect 110708 16546 111012 16574
rect 110512 8968 110564 8974
rect 110512 8910 110564 8916
rect 110432 6886 110552 6914
rect 109684 3664 109736 3670
rect 109684 3606 109736 3612
rect 108304 3596 108356 3602
rect 108304 3538 108356 3544
rect 109316 3596 109368 3602
rect 109316 3538 109368 3544
rect 106832 3460 106884 3466
rect 106832 3402 106884 3408
rect 106936 480 106964 3470
rect 107672 3454 108160 3482
rect 108132 480 108160 3454
rect 109328 480 109356 3538
rect 110524 480 110552 6886
rect 110984 3482 111012 16546
rect 111076 3602 111104 78066
rect 111444 77178 111472 79750
rect 111812 77994 111840 79886
rect 111984 79824 112036 79830
rect 112226 79778 112254 80036
rect 112594 79830 112622 80036
rect 111984 79766 112036 79772
rect 111800 77988 111852 77994
rect 111800 77930 111852 77936
rect 111892 77308 111944 77314
rect 111892 77250 111944 77256
rect 111432 77172 111484 77178
rect 111432 77114 111484 77120
rect 111064 3596 111116 3602
rect 111064 3538 111116 3544
rect 111904 3534 111932 77250
rect 111996 4214 112024 79766
rect 112088 79750 112254 79778
rect 112582 79824 112634 79830
rect 112962 79778 112990 80036
rect 113330 79914 113358 80036
rect 113698 79914 113726 80036
rect 114066 79914 114094 80036
rect 112582 79766 112634 79772
rect 112916 79750 112990 79778
rect 113284 79886 113358 79914
rect 113652 79886 113726 79914
rect 114020 79886 114094 79914
rect 112088 22166 112116 79750
rect 112168 78668 112220 78674
rect 112168 78610 112220 78616
rect 112076 22160 112128 22166
rect 112076 22102 112128 22108
rect 112180 16574 112208 78610
rect 112916 77314 112944 79750
rect 113284 77858 113312 79886
rect 113652 78130 113680 79886
rect 114020 78402 114048 79886
rect 114434 79778 114462 80036
rect 114802 79914 114830 80036
rect 114388 79750 114462 79778
rect 114572 79886 114830 79914
rect 114008 78396 114060 78402
rect 114008 78338 114060 78344
rect 113640 78124 113692 78130
rect 113640 78066 113692 78072
rect 113272 77852 113324 77858
rect 113272 77794 113324 77800
rect 112904 77308 112956 77314
rect 112904 77250 112956 77256
rect 114388 60734 114416 79750
rect 114572 78674 114600 79886
rect 115170 79778 115198 80036
rect 115538 79778 115566 80036
rect 114664 79750 115198 79778
rect 115492 79750 115566 79778
rect 115912 79778 115940 80036
rect 116032 79824 116084 79830
rect 115912 79750 115980 79778
rect 116182 79778 116210 80036
rect 116550 79778 116578 80036
rect 116918 79830 116946 80036
rect 116032 79766 116084 79772
rect 114560 78668 114612 78674
rect 114560 78610 114612 78616
rect 113376 60706 114416 60734
rect 113376 23458 113404 60706
rect 113364 23452 113416 23458
rect 113364 23394 113416 23400
rect 112180 16546 112392 16574
rect 111984 4208 112036 4214
rect 111984 4150 112036 4156
rect 111892 3528 111944 3534
rect 110984 3454 111656 3482
rect 111892 3470 111944 3476
rect 111628 480 111656 3454
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114664 6914 114692 79750
rect 115492 60734 115520 79750
rect 114572 6886 114692 6914
rect 114756 60706 115520 60734
rect 114572 2802 114600 6886
rect 114480 2774 114600 2802
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 354 114090 480
rect 114480 354 114508 2774
rect 113978 326 114508 354
rect 114756 354 114784 60706
rect 115952 3346 115980 79750
rect 116044 3466 116072 79766
rect 116136 79750 116210 79778
rect 116320 79750 116578 79778
rect 116906 79824 116958 79830
rect 116906 79766 116958 79772
rect 117292 79778 117320 80036
rect 117654 79778 117682 80036
rect 117292 79750 117360 79778
rect 116136 3534 116164 79750
rect 116320 60734 116348 79750
rect 117332 74610 117360 79750
rect 117608 79750 117682 79778
rect 118028 79778 118056 80036
rect 118396 79778 118424 80036
rect 118758 79778 118786 80036
rect 119494 79778 119522 80036
rect 119862 79778 119890 80036
rect 118028 79750 118096 79778
rect 118396 79750 118464 79778
rect 117332 74582 117452 74610
rect 117424 67634 117452 74582
rect 117608 74534 117636 79750
rect 118068 77382 118096 79750
rect 118436 77790 118464 79750
rect 118712 79750 118786 79778
rect 118896 79750 119522 79778
rect 119816 79750 119890 79778
rect 120604 79778 120632 80036
rect 120972 79778 121000 80036
rect 121340 79778 121368 80036
rect 121552 79892 121604 79898
rect 121552 79834 121604 79840
rect 121460 79824 121512 79830
rect 120604 79750 120672 79778
rect 120972 79750 121040 79778
rect 121340 79750 121408 79778
rect 121460 79766 121512 79772
rect 118424 77784 118476 77790
rect 118424 77726 118476 77732
rect 118056 77376 118108 77382
rect 118056 77318 118108 77324
rect 117332 67606 117452 67634
rect 117516 74506 117636 74534
rect 117332 62914 117360 67606
rect 117332 62886 117452 62914
rect 117320 62824 117372 62830
rect 117320 62766 117372 62772
rect 116228 60706 116348 60734
rect 116228 9654 116256 60706
rect 116216 9648 116268 9654
rect 116216 9590 116268 9596
rect 117332 8294 117360 62766
rect 117424 11014 117452 62886
rect 117516 62830 117544 74506
rect 117504 62824 117556 62830
rect 117504 62766 117556 62772
rect 117412 11008 117464 11014
rect 117412 10950 117464 10956
rect 117320 8288 117372 8294
rect 117320 8230 117372 8236
rect 118712 4962 118740 79750
rect 118792 77308 118844 77314
rect 118792 77250 118844 77256
rect 118804 12866 118832 77250
rect 118896 13122 118924 79750
rect 119344 77376 119396 77382
rect 119344 77318 119396 77324
rect 118884 13116 118936 13122
rect 118884 13058 118936 13064
rect 118804 12838 118924 12866
rect 118792 9648 118844 9654
rect 118792 9590 118844 9596
rect 118700 4956 118752 4962
rect 118700 4898 118752 4904
rect 116124 3528 116176 3534
rect 116124 3470 116176 3476
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 116032 3460 116084 3466
rect 116032 3402 116084 3408
rect 115952 3318 116440 3346
rect 116412 480 116440 3318
rect 117608 480 117636 3470
rect 118804 480 118832 9590
rect 118896 9178 118924 12838
rect 118884 9172 118936 9178
rect 118884 9114 118936 9120
rect 119356 4146 119384 77318
rect 119816 77314 119844 79750
rect 120644 78062 120672 79750
rect 120632 78056 120684 78062
rect 120632 77998 120684 78004
rect 121012 77314 121040 79750
rect 121380 77858 121408 79750
rect 121368 77852 121420 77858
rect 121368 77794 121420 77800
rect 119804 77308 119856 77314
rect 119804 77250 119856 77256
rect 121000 77308 121052 77314
rect 121000 77250 121052 77256
rect 120632 11008 120684 11014
rect 120632 10950 120684 10956
rect 119344 4140 119396 4146
rect 119344 4082 119396 4088
rect 119896 3460 119948 3466
rect 119896 3402 119948 3408
rect 119908 480 119936 3402
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 113978 -960 114090 326
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 10950
rect 121472 4894 121500 79766
rect 121564 7818 121592 79834
rect 121702 79778 121730 80036
rect 122070 79830 122098 80036
rect 122438 79898 122466 80036
rect 122426 79892 122478 79898
rect 122426 79834 122478 79840
rect 121656 79750 121730 79778
rect 122058 79824 122110 79830
rect 122812 79812 122840 80036
rect 122812 79784 122972 79812
rect 122058 79766 122110 79772
rect 121552 7812 121604 7818
rect 121552 7754 121604 7760
rect 121656 7682 121684 79750
rect 122840 79688 122892 79694
rect 122840 79630 122892 79636
rect 122104 77308 122156 77314
rect 122104 77250 122156 77256
rect 122116 8974 122144 77250
rect 122852 10402 122880 79630
rect 122944 15910 122972 79784
rect 123180 79642 123208 80036
rect 123542 79898 123570 80036
rect 123530 79892 123582 79898
rect 123530 79834 123582 79840
rect 123910 79778 123938 80036
rect 124278 79914 124306 80036
rect 123312 79750 123938 79778
rect 124232 79886 124306 79914
rect 123180 79614 123248 79642
rect 123220 77382 123248 79614
rect 123208 77376 123260 77382
rect 123208 77318 123260 77324
rect 123312 64874 123340 79750
rect 124232 77926 124260 79886
rect 124312 79824 124364 79830
rect 124646 79778 124674 80036
rect 125014 79778 125042 80036
rect 125382 79830 125410 80036
rect 124312 79766 124364 79772
rect 124220 77920 124272 77926
rect 124220 77862 124272 77868
rect 123484 77852 123536 77858
rect 123484 77794 123536 77800
rect 123036 64846 123340 64874
rect 123036 17474 123064 64846
rect 123024 17468 123076 17474
rect 123024 17410 123076 17416
rect 122932 15904 122984 15910
rect 122932 15846 122984 15852
rect 122840 10396 122892 10402
rect 122840 10338 122892 10344
rect 123496 9042 123524 77794
rect 124220 77784 124272 77790
rect 124220 77726 124272 77732
rect 123484 9036 123536 9042
rect 123484 8978 123536 8984
rect 122104 8968 122156 8974
rect 122104 8910 122156 8916
rect 122288 8288 122340 8294
rect 122288 8230 122340 8236
rect 121644 7676 121696 7682
rect 121644 7618 121696 7624
rect 121460 4888 121512 4894
rect 121460 4830 121512 4836
rect 122300 480 122328 8230
rect 123484 4140 123536 4146
rect 123484 4082 123536 4088
rect 123496 480 123524 4082
rect 124232 1306 124260 77726
rect 124324 4826 124352 79766
rect 124416 79750 124674 79778
rect 124968 79750 125042 79778
rect 125370 79824 125422 79830
rect 125750 79778 125778 80036
rect 126118 79778 126146 80036
rect 126486 79778 126514 80036
rect 126854 79778 126882 80036
rect 125370 79766 125422 79772
rect 125612 79750 125778 79778
rect 125888 79750 126146 79778
rect 126440 79750 126514 79778
rect 126808 79750 126882 79778
rect 126980 79824 127032 79830
rect 127222 79778 127250 80036
rect 127590 79778 127618 80036
rect 126980 79766 127032 79772
rect 124416 9110 124444 79750
rect 124968 64874 124996 79750
rect 124508 64846 124996 64874
rect 124508 18630 124536 64846
rect 124496 18624 124548 18630
rect 124496 18566 124548 18572
rect 125612 10334 125640 79750
rect 125784 77308 125836 77314
rect 125784 77250 125836 77256
rect 125692 77240 125744 77246
rect 125692 77182 125744 77188
rect 125704 11762 125732 77182
rect 125796 11898 125824 77250
rect 125888 42090 125916 79750
rect 126244 78056 126296 78062
rect 126244 77998 126296 78004
rect 125876 42084 125928 42090
rect 125876 42026 125928 42032
rect 125784 11892 125836 11898
rect 125784 11834 125836 11840
rect 125692 11756 125744 11762
rect 125692 11698 125744 11704
rect 125600 10328 125652 10334
rect 125600 10270 125652 10276
rect 124404 9104 124456 9110
rect 124404 9046 124456 9052
rect 126256 5574 126284 77998
rect 126440 77314 126468 79750
rect 126428 77308 126480 77314
rect 126428 77250 126480 77256
rect 126808 77246 126836 79750
rect 126796 77240 126848 77246
rect 126796 77182 126848 77188
rect 126992 6322 127020 79766
rect 127084 79750 127250 79778
rect 127544 79750 127618 79778
rect 127964 79778 127992 80036
rect 128234 79830 128262 80036
rect 128222 79824 128274 79830
rect 127964 79750 128032 79778
rect 128602 79778 128630 80036
rect 128970 79778 128998 80036
rect 128222 79766 128274 79772
rect 126980 6316 127032 6322
rect 126980 6258 127032 6264
rect 126980 6180 127032 6186
rect 126980 6122 127032 6128
rect 126244 5568 126296 5574
rect 126244 5510 126296 5516
rect 125876 4956 125928 4962
rect 125876 4898 125928 4904
rect 124312 4820 124364 4826
rect 124312 4762 124364 4768
rect 124232 1278 124720 1306
rect 124692 480 124720 1278
rect 125888 480 125916 4898
rect 126992 480 127020 6122
rect 127084 5982 127112 79750
rect 127544 64874 127572 79750
rect 128004 77314 128032 79750
rect 128372 79750 128630 79778
rect 128740 79750 128998 79778
rect 129344 79778 129372 80036
rect 129712 79778 129740 80036
rect 129924 79824 129976 79830
rect 129344 79750 129412 79778
rect 129712 79750 129872 79778
rect 130074 79778 130102 80036
rect 130442 79778 130470 80036
rect 130810 79830 130838 80036
rect 129924 79766 129976 79772
rect 127992 77308 128044 77314
rect 127992 77250 128044 77256
rect 127176 64846 127572 64874
rect 127176 11830 127204 64846
rect 128372 13258 128400 79750
rect 128740 64874 128768 79750
rect 129384 78130 129412 79750
rect 129372 78124 129424 78130
rect 129372 78066 129424 78072
rect 129096 77920 129148 77926
rect 129096 77862 129148 77868
rect 129004 77376 129056 77382
rect 129004 77318 129056 77324
rect 128464 64846 128768 64874
rect 128360 13252 128412 13258
rect 128360 13194 128412 13200
rect 128464 13190 128492 64846
rect 128452 13184 128504 13190
rect 128452 13126 128504 13132
rect 128176 13116 128228 13122
rect 128176 13058 128228 13064
rect 127164 11824 127216 11830
rect 127164 11766 127216 11772
rect 127164 6316 127216 6322
rect 127164 6258 127216 6264
rect 127072 5976 127124 5982
rect 127072 5918 127124 5924
rect 127176 3466 127204 6258
rect 127164 3460 127216 3466
rect 127164 3402 127216 3408
rect 128188 480 128216 13058
rect 128360 5976 128412 5982
rect 128360 5918 128412 5924
rect 128372 3602 128400 5918
rect 129016 4962 129044 77318
rect 129108 10470 129136 77862
rect 129188 77308 129240 77314
rect 129188 77250 129240 77256
rect 129740 77308 129792 77314
rect 129740 77250 129792 77256
rect 129200 40866 129228 77250
rect 129188 40860 129240 40866
rect 129188 40802 129240 40808
rect 129752 13122 129780 77250
rect 129844 14618 129872 79750
rect 129832 14612 129884 14618
rect 129832 14554 129884 14560
rect 129936 14550 129964 79766
rect 130028 79750 130102 79778
rect 130396 79750 130470 79778
rect 130798 79824 130850 79830
rect 131178 79778 131206 80036
rect 131552 79880 131580 80036
rect 131920 79880 131948 80036
rect 131552 79852 131620 79880
rect 131920 79852 131988 79880
rect 130798 79766 130850 79772
rect 131132 79750 131206 79778
rect 130028 19990 130056 79750
rect 130396 77314 130424 79750
rect 130384 77308 130436 77314
rect 130384 77250 130436 77256
rect 130016 19984 130068 19990
rect 130016 19926 130068 19932
rect 129924 14544 129976 14550
rect 129924 14486 129976 14492
rect 129740 13116 129792 13122
rect 129740 13058 129792 13064
rect 129096 10464 129148 10470
rect 129096 10406 129148 10412
rect 129372 9172 129424 9178
rect 129372 9114 129424 9120
rect 129004 4956 129056 4962
rect 129004 4898 129056 4904
rect 128360 3596 128412 3602
rect 128360 3538 128412 3544
rect 129384 480 129412 9114
rect 130568 7608 130620 7614
rect 130568 7550 130620 7556
rect 130580 480 130608 7550
rect 131132 6254 131160 79750
rect 131592 78538 131620 79852
rect 131580 78532 131632 78538
rect 131580 78474 131632 78480
rect 131960 77994 131988 79852
rect 132282 79778 132310 80036
rect 132236 79750 132310 79778
rect 132500 79824 132552 79830
rect 132500 79766 132552 79772
rect 132656 79778 132684 80036
rect 133018 79830 133046 80036
rect 133006 79824 133058 79830
rect 131948 77988 132000 77994
rect 131948 77930 132000 77936
rect 132236 64874 132264 79750
rect 131224 64846 132264 64874
rect 131224 6390 131252 64846
rect 132512 14482 132540 79766
rect 132656 79750 132816 79778
rect 133386 79778 133414 80036
rect 133754 79778 133782 80036
rect 134122 79914 134150 80036
rect 133006 79766 133058 79772
rect 132684 77308 132736 77314
rect 132684 77250 132736 77256
rect 132592 77240 132644 77246
rect 132592 77182 132644 77188
rect 132604 20058 132632 77182
rect 132696 21486 132724 77250
rect 132788 27062 132816 79750
rect 133340 79750 133414 79778
rect 133708 79750 133782 79778
rect 133892 79886 134150 79914
rect 133340 77314 133368 79750
rect 133328 77308 133380 77314
rect 133328 77250 133380 77256
rect 133708 77246 133736 79750
rect 133696 77240 133748 77246
rect 133696 77182 133748 77188
rect 132776 27056 132828 27062
rect 132776 26998 132828 27004
rect 132684 21480 132736 21486
rect 132684 21422 132736 21428
rect 132592 20052 132644 20058
rect 132592 19994 132644 20000
rect 133892 15978 133920 79886
rect 133972 79824 134024 79830
rect 134490 79778 134518 80036
rect 134858 79830 134886 80036
rect 135232 79914 135260 80036
rect 135600 79914 135628 80036
rect 135232 79886 135392 79914
rect 135600 79886 135668 79914
rect 133972 79766 134024 79772
rect 133984 20126 134012 79766
rect 134076 79750 134518 79778
rect 134846 79824 134898 79830
rect 134846 79766 134898 79772
rect 134076 21418 134104 79750
rect 134524 78532 134576 78538
rect 134524 78474 134576 78480
rect 134536 24206 134564 78474
rect 135364 77382 135392 79886
rect 135640 77450 135668 79886
rect 135962 79778 135990 80036
rect 135732 79750 135990 79778
rect 136336 79778 136364 80036
rect 136704 79778 136732 80036
rect 137066 79778 137094 80036
rect 137434 79778 137462 80036
rect 137802 79778 137830 80036
rect 138170 79778 138198 80036
rect 138538 79778 138566 80036
rect 138906 79778 138934 80036
rect 139274 79778 139302 80036
rect 139642 79914 139670 80036
rect 136336 79750 136404 79778
rect 136704 79750 136864 79778
rect 135628 77444 135680 77450
rect 135628 77386 135680 77392
rect 135352 77376 135404 77382
rect 135352 77318 135404 77324
rect 135732 64874 135760 79750
rect 136376 78198 136404 79750
rect 136364 78192 136416 78198
rect 136364 78134 136416 78140
rect 135904 78124 135956 78130
rect 135904 78066 135956 78072
rect 135272 64846 135760 64874
rect 135272 40798 135300 64846
rect 135260 40792 135312 40798
rect 135260 40734 135312 40740
rect 134524 24200 134576 24206
rect 134524 24142 134576 24148
rect 134064 21412 134116 21418
rect 134064 21354 134116 21360
rect 133972 20120 134024 20126
rect 133972 20062 134024 20068
rect 133880 15972 133932 15978
rect 133880 15914 133932 15920
rect 132500 14476 132552 14482
rect 132500 14418 132552 14424
rect 134156 9036 134208 9042
rect 134156 8978 134208 8984
rect 132960 8968 133012 8974
rect 132960 8910 133012 8916
rect 131212 6384 131264 6390
rect 131212 6326 131264 6332
rect 131120 6248 131172 6254
rect 131120 6190 131172 6196
rect 131764 5568 131816 5574
rect 131764 5510 131816 5516
rect 131776 480 131804 5510
rect 132972 480 133000 8910
rect 134168 480 134196 8978
rect 135260 7676 135312 7682
rect 135260 7618 135312 7624
rect 135272 480 135300 7618
rect 135916 3534 135944 78066
rect 136732 77308 136784 77314
rect 136732 77250 136784 77256
rect 136640 77240 136692 77246
rect 136640 77182 136692 77188
rect 136652 7682 136680 77182
rect 136744 16046 136772 77250
rect 136836 24138 136864 79750
rect 136928 79750 137094 79778
rect 137388 79750 137462 79778
rect 137756 79750 137830 79778
rect 138032 79750 138198 79778
rect 138308 79750 138566 79778
rect 138860 79750 138934 79778
rect 139228 79750 139302 79778
rect 139412 79886 139670 79914
rect 140010 79898 140038 80036
rect 139998 79892 140050 79898
rect 136928 28354 136956 79750
rect 137284 77376 137336 77382
rect 137284 77318 137336 77324
rect 137296 50386 137324 77318
rect 137388 77314 137416 79750
rect 137376 77308 137428 77314
rect 137376 77250 137428 77256
rect 137756 77246 137784 79750
rect 137744 77240 137796 77246
rect 137744 77182 137796 77188
rect 137284 50380 137336 50386
rect 137284 50322 137336 50328
rect 136916 28348 136968 28354
rect 136916 28290 136968 28296
rect 136824 24132 136876 24138
rect 136824 24074 136876 24080
rect 136732 16040 136784 16046
rect 136732 15982 136784 15988
rect 137652 7812 137704 7818
rect 137652 7754 137704 7760
rect 136640 7676 136692 7682
rect 136640 7618 136692 7624
rect 136456 4888 136508 4894
rect 136456 4830 136508 4836
rect 135904 3528 135956 3534
rect 135904 3470 135956 3476
rect 136468 480 136496 4830
rect 137664 480 137692 7754
rect 138032 7750 138060 79750
rect 138204 77308 138256 77314
rect 138204 77250 138256 77256
rect 138112 77240 138164 77246
rect 138112 77182 138164 77188
rect 138124 25566 138152 77182
rect 138216 29782 138244 77250
rect 138308 44946 138336 79750
rect 138860 77246 138888 79750
rect 139228 77314 139256 79750
rect 139216 77308 139268 77314
rect 139216 77250 139268 77256
rect 138848 77240 138900 77246
rect 138848 77182 138900 77188
rect 138296 44940 138348 44946
rect 138296 44882 138348 44888
rect 138204 29776 138256 29782
rect 138204 29718 138256 29724
rect 138112 25560 138164 25566
rect 138112 25502 138164 25508
rect 139412 15910 139440 79886
rect 139998 79834 140050 79840
rect 139584 79824 139636 79830
rect 140286 79778 140314 80036
rect 140654 79778 140682 80036
rect 139584 79766 139636 79772
rect 139492 77308 139544 77314
rect 139492 77250 139544 77256
rect 139504 17406 139532 77250
rect 139596 26994 139624 79766
rect 139688 79750 140314 79778
rect 140608 79750 140682 79778
rect 140780 79824 140832 79830
rect 141022 79778 141050 80036
rect 141390 79778 141418 80036
rect 141758 79830 141786 80036
rect 140780 79766 140832 79772
rect 139688 31142 139716 79750
rect 140608 77314 140636 79750
rect 140596 77308 140648 77314
rect 140596 77250 140648 77256
rect 139676 31136 139728 31142
rect 139676 31078 139728 31084
rect 139584 26988 139636 26994
rect 139584 26930 139636 26936
rect 139492 17400 139544 17406
rect 139492 17342 139544 17348
rect 140792 17338 140820 79766
rect 140884 79750 141050 79778
rect 141160 79750 141418 79778
rect 141746 79824 141798 79830
rect 142132 79812 142160 80036
rect 142132 79784 142384 79812
rect 141746 79766 141798 79772
rect 140884 28286 140912 79750
rect 141160 64874 141188 79750
rect 141424 77988 141476 77994
rect 141424 77930 141476 77936
rect 140976 64846 141188 64874
rect 140976 35358 141004 64846
rect 140964 35352 141016 35358
rect 140964 35294 141016 35300
rect 140872 28280 140924 28286
rect 140872 28222 140924 28228
rect 141436 22778 141464 77930
rect 142356 77738 142384 79784
rect 142500 79778 142528 80036
rect 142862 79778 142890 80036
rect 143230 79778 143258 80036
rect 143598 79778 143626 80036
rect 143972 79880 144000 80036
rect 143972 79852 144040 79880
rect 142500 79750 142568 79778
rect 142356 77710 142476 77738
rect 142158 77480 142214 77489
rect 142448 77450 142476 77710
rect 142540 77489 142568 79750
rect 142632 79750 142890 79778
rect 143000 79750 143258 79778
rect 143552 79750 143626 79778
rect 142526 77480 142582 77489
rect 142158 77415 142214 77424
rect 142436 77444 142488 77450
rect 141424 22772 141476 22778
rect 141424 22714 141476 22720
rect 140780 17332 140832 17338
rect 140780 17274 140832 17280
rect 138848 15904 138900 15910
rect 138848 15846 138900 15852
rect 139400 15904 139452 15910
rect 139400 15846 139452 15852
rect 138020 7744 138072 7750
rect 138020 7686 138072 7692
rect 138860 480 138888 15846
rect 141240 10396 141292 10402
rect 141240 10338 141292 10344
rect 140044 4956 140096 4962
rect 140044 4898 140096 4904
rect 140056 480 140084 4898
rect 141252 480 141280 10338
rect 142172 9042 142200 77415
rect 142526 77415 142582 77424
rect 142436 77386 142488 77392
rect 142632 77330 142660 79750
rect 142264 77302 142660 77330
rect 142264 17270 142292 77302
rect 143000 77194 143028 79750
rect 142356 77166 143028 77194
rect 142356 29646 142384 77166
rect 142436 77104 142488 77110
rect 142436 77046 142488 77052
rect 142448 29714 142476 77046
rect 142436 29708 142488 29714
rect 142436 29650 142488 29656
rect 142344 29640 142396 29646
rect 142344 29582 142396 29588
rect 142344 17468 142396 17474
rect 142344 17410 142396 17416
rect 142252 17264 142304 17270
rect 142252 17206 142304 17212
rect 142356 16574 142384 17410
rect 142356 16546 142476 16574
rect 142160 9036 142212 9042
rect 142160 8978 142212 8984
rect 142448 480 142476 16546
rect 143552 12782 143580 79750
rect 144012 77994 144040 79852
rect 144334 79778 144362 80036
rect 144702 79778 144730 80036
rect 144104 79750 144362 79778
rect 144656 79750 144730 79778
rect 144920 79824 144972 79830
rect 145070 79778 145098 80036
rect 145438 79778 145466 80036
rect 145806 79778 145834 80036
rect 146174 79830 146202 80036
rect 146300 79892 146352 79898
rect 146300 79834 146352 79840
rect 144920 79766 144972 79772
rect 144000 77988 144052 77994
rect 144000 77930 144052 77936
rect 143632 77308 143684 77314
rect 143632 77250 143684 77256
rect 143540 12776 143592 12782
rect 143540 12718 143592 12724
rect 143540 10464 143592 10470
rect 143540 10406 143592 10412
rect 143552 480 143580 10406
rect 143644 9314 143672 77250
rect 144104 64874 144132 79750
rect 144184 77512 144236 77518
rect 144184 77454 144236 77460
rect 143736 64846 144132 64874
rect 143736 31074 143764 64846
rect 143724 31068 143776 31074
rect 143724 31010 143776 31016
rect 144196 21554 144224 77454
rect 144656 77314 144684 79750
rect 144644 77308 144696 77314
rect 144644 77250 144696 77256
rect 144184 21548 144236 21554
rect 144184 21490 144236 21496
rect 144932 18766 144960 79766
rect 145024 79750 145098 79778
rect 145208 79750 145466 79778
rect 145760 79750 145834 79778
rect 146162 79824 146214 79830
rect 146162 79766 146214 79772
rect 145024 40730 145052 79750
rect 145104 77308 145156 77314
rect 145104 77250 145156 77256
rect 145116 43450 145144 77250
rect 145208 44878 145236 79750
rect 145760 77314 145788 79750
rect 145748 77308 145800 77314
rect 145748 77250 145800 77256
rect 145196 44872 145248 44878
rect 145196 44814 145248 44820
rect 145104 43444 145156 43450
rect 145104 43386 145156 43392
rect 145012 40724 145064 40730
rect 145012 40666 145064 40672
rect 144920 18760 144972 18766
rect 144920 18702 144972 18708
rect 144920 18624 144972 18630
rect 144920 18566 144972 18572
rect 144932 16574 144960 18566
rect 144932 16546 145512 16574
rect 143724 12776 143776 12782
rect 143724 12718 143776 12724
rect 143632 9308 143684 9314
rect 143632 9250 143684 9256
rect 143736 8974 143764 12718
rect 144736 9104 144788 9110
rect 144736 9046 144788 9052
rect 143724 8968 143776 8974
rect 143724 8910 143776 8916
rect 144748 480 144776 9046
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 146312 4962 146340 79834
rect 146392 79824 146444 79830
rect 146542 79778 146570 80036
rect 146910 79830 146938 80036
rect 147278 79898 147306 80036
rect 147266 79892 147318 79898
rect 147266 79834 147318 79840
rect 146392 79766 146444 79772
rect 146404 10402 146432 79766
rect 146496 79750 146570 79778
rect 146898 79824 146950 79830
rect 146898 79766 146950 79772
rect 147652 79778 147680 80036
rect 147864 79824 147916 79830
rect 147652 79750 147812 79778
rect 148014 79778 148042 80036
rect 148382 79778 148410 80036
rect 148750 79830 148778 80036
rect 147864 79766 147916 79772
rect 146496 32434 146524 79750
rect 147680 77308 147732 77314
rect 147680 77250 147732 77256
rect 146484 32428 146536 32434
rect 146484 32370 146536 32376
rect 146392 10396 146444 10402
rect 146392 10338 146444 10344
rect 146300 4956 146352 4962
rect 146300 4898 146352 4904
rect 147692 4894 147720 77250
rect 147784 33794 147812 79750
rect 147876 35290 147904 79766
rect 147968 79750 148042 79778
rect 148336 79750 148410 79778
rect 148738 79824 148790 79830
rect 148738 79766 148790 79772
rect 149124 79778 149152 80036
rect 149492 79880 149520 80036
rect 149492 79852 149560 79880
rect 149124 79750 149192 79778
rect 147968 47598 147996 79750
rect 148336 77314 148364 79750
rect 148324 77308 148376 77314
rect 148324 77250 148376 77256
rect 149060 77308 149112 77314
rect 149060 77250 149112 77256
rect 147956 47592 148008 47598
rect 147956 47534 148008 47540
rect 147864 35284 147916 35290
rect 147864 35226 147916 35232
rect 147772 33788 147824 33794
rect 147772 33730 147824 33736
rect 149072 10334 149100 77250
rect 149164 60042 149192 79750
rect 149532 78062 149560 79852
rect 149854 79778 149882 80036
rect 150222 79778 150250 80036
rect 150590 79778 150618 80036
rect 150958 79778 150986 80036
rect 151326 79778 151354 80036
rect 151694 79778 151722 80036
rect 152062 79914 152090 80036
rect 151820 79892 151872 79898
rect 151820 79834 151872 79840
rect 151924 79886 152090 79914
rect 149716 79750 149882 79778
rect 150176 79750 150250 79778
rect 150452 79750 150618 79778
rect 150728 79750 150986 79778
rect 151280 79750 151354 79778
rect 151648 79750 151722 79778
rect 149520 78056 149572 78062
rect 149520 77998 149572 78004
rect 149716 64874 149744 79750
rect 150176 77314 150204 79750
rect 150164 77308 150216 77314
rect 150164 77250 150216 77256
rect 149256 64846 149744 64874
rect 149152 60036 149204 60042
rect 149152 59978 149204 59984
rect 149256 42090 149284 64846
rect 149152 42084 149204 42090
rect 149152 42026 149204 42032
rect 149244 42084 149296 42090
rect 149244 42026 149296 42032
rect 149164 16574 149192 42026
rect 149164 16546 149560 16574
rect 147864 10328 147916 10334
rect 147864 10270 147916 10276
rect 149060 10328 149112 10334
rect 149060 10270 149112 10276
rect 147680 4888 147732 4894
rect 147680 4830 147732 4836
rect 147128 4820 147180 4826
rect 147128 4762 147180 4768
rect 147140 480 147168 4762
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 10270
rect 149532 480 149560 16546
rect 150452 4826 150480 79750
rect 150624 77308 150676 77314
rect 150624 77250 150676 77256
rect 150532 77240 150584 77246
rect 150532 77182 150584 77188
rect 150544 10674 150572 77182
rect 150636 18698 150664 77250
rect 150728 26926 150756 79750
rect 151280 77246 151308 79750
rect 151648 77314 151676 79750
rect 151636 77308 151688 77314
rect 151636 77250 151688 77256
rect 151268 77240 151320 77246
rect 151268 77182 151320 77188
rect 150716 26920 150768 26926
rect 150716 26862 150768 26868
rect 150624 18692 150676 18698
rect 150624 18634 150676 18640
rect 151832 18630 151860 79834
rect 151924 35222 151952 79886
rect 152004 79824 152056 79830
rect 152338 79778 152366 80036
rect 152706 79898 152734 80036
rect 152694 79892 152746 79898
rect 152694 79834 152746 79840
rect 153074 79830 153102 80036
rect 152004 79766 152056 79772
rect 152016 36922 152044 79766
rect 152108 79750 152366 79778
rect 153062 79824 153114 79830
rect 153062 79766 153114 79772
rect 153200 79824 153252 79830
rect 153442 79778 153470 80036
rect 153200 79766 153252 79772
rect 152108 50726 152136 79750
rect 152096 50720 152148 50726
rect 152096 50662 152148 50668
rect 153212 38282 153240 79766
rect 153304 79750 153470 79778
rect 153816 79778 153844 80036
rect 154178 79830 154206 80036
rect 154166 79824 154218 79830
rect 153816 79750 153884 79778
rect 154166 79766 154218 79772
rect 154552 79778 154580 80036
rect 154914 79778 154942 80036
rect 155282 79778 155310 80036
rect 155650 79778 155678 80036
rect 154552 79750 154712 79778
rect 153304 52086 153332 79750
rect 153856 78130 153884 79750
rect 153844 78124 153896 78130
rect 153844 78066 153896 78072
rect 154580 77308 154632 77314
rect 154580 77250 154632 77256
rect 153292 52080 153344 52086
rect 153292 52022 153344 52028
rect 153200 38276 153252 38282
rect 153200 38218 153252 38224
rect 152004 36916 152056 36922
rect 152004 36858 152056 36864
rect 151912 35216 151964 35222
rect 151912 35158 151964 35164
rect 151820 18624 151872 18630
rect 151820 18566 151872 18572
rect 150624 11892 150676 11898
rect 150624 11834 150676 11840
rect 150532 10668 150584 10674
rect 150532 10610 150584 10616
rect 150440 4820 150492 4826
rect 150440 4762 150492 4768
rect 150636 480 150664 11834
rect 154592 11830 154620 77250
rect 154684 11898 154712 79750
rect 154776 79750 154942 79778
rect 155052 79750 155310 79778
rect 155604 79750 155678 79778
rect 156024 79778 156052 80036
rect 156144 79824 156196 79830
rect 156024 79750 156092 79778
rect 156386 79778 156414 80036
rect 156754 79778 156782 80036
rect 157122 79830 157150 80036
rect 157340 79892 157392 79898
rect 157340 79834 157392 79840
rect 156144 79766 156196 79772
rect 154776 24546 154804 79750
rect 155052 64874 155080 79750
rect 155604 77314 155632 79750
rect 155592 77308 155644 77314
rect 155592 77250 155644 77256
rect 155960 77308 156012 77314
rect 155960 77250 156012 77256
rect 154960 64846 155080 64874
rect 154856 40860 154908 40866
rect 154856 40802 154908 40808
rect 154764 24540 154816 24546
rect 154764 24482 154816 24488
rect 154868 16574 154896 40802
rect 154960 39370 154988 64846
rect 154948 39364 155000 39370
rect 154948 39306 155000 39312
rect 154868 16546 155448 16574
rect 154672 11892 154724 11898
rect 154672 11834 154724 11840
rect 153752 11824 153804 11830
rect 153752 11766 153804 11772
rect 154580 11824 154632 11830
rect 154580 11766 154632 11772
rect 151820 11756 151872 11762
rect 151820 11698 151872 11704
rect 151832 480 151860 11698
rect 153016 3596 153068 3602
rect 153016 3538 153068 3544
rect 153028 480 153056 3538
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 11766
rect 155420 480 155448 16546
rect 155972 11762 156000 77250
rect 156064 24478 156092 79750
rect 156156 25906 156184 79766
rect 156248 79750 156414 79778
rect 156708 79750 156782 79778
rect 157110 79824 157162 79830
rect 157110 79766 157162 79772
rect 156248 43790 156276 79750
rect 156708 77314 156736 79750
rect 156696 77308 156748 77314
rect 156696 77250 156748 77256
rect 156236 43784 156288 43790
rect 156236 43726 156288 43732
rect 156144 25900 156196 25906
rect 156144 25842 156196 25848
rect 156052 24472 156104 24478
rect 156052 24414 156104 24420
rect 157352 13462 157380 79834
rect 157496 79778 157524 80036
rect 157858 79898 157886 80036
rect 158226 79898 158254 80036
rect 157846 79892 157898 79898
rect 157846 79834 157898 79840
rect 158214 79892 158266 79898
rect 158214 79834 158266 79840
rect 158594 79778 158622 80036
rect 158962 79778 158990 80036
rect 159330 79778 159358 80036
rect 159698 79778 159726 80036
rect 157496 79750 157564 79778
rect 157432 79688 157484 79694
rect 157432 79630 157484 79636
rect 157444 25838 157472 79630
rect 157536 46510 157564 79750
rect 157628 79750 158622 79778
rect 158732 79750 158990 79778
rect 159100 79750 159358 79778
rect 159468 79750 159726 79778
rect 160072 79778 160100 80036
rect 160434 79778 160462 80036
rect 160802 79778 160830 80036
rect 161170 79778 161198 80036
rect 161538 79778 161566 80036
rect 161906 79778 161934 80036
rect 162274 79778 162302 80036
rect 162642 79778 162670 80036
rect 160072 79750 160140 79778
rect 157628 47938 157656 79750
rect 157616 47932 157668 47938
rect 157616 47874 157668 47880
rect 157524 46504 157576 46510
rect 157524 46446 157576 46452
rect 157432 25832 157484 25838
rect 157432 25774 157484 25780
rect 157340 13456 157392 13462
rect 157340 13398 157392 13404
rect 158732 13326 158760 79750
rect 159100 70394 159128 79750
rect 158824 70366 159128 70394
rect 158824 22982 158852 70366
rect 159468 64874 159496 79750
rect 160112 75426 160140 79750
rect 160020 75398 160140 75426
rect 160204 79750 160462 79778
rect 160756 79750 160830 79778
rect 160940 79750 161198 79778
rect 161492 79750 161566 79778
rect 161676 79750 161934 79778
rect 162044 79750 162302 79778
rect 162596 79750 162670 79778
rect 162860 79824 162912 79830
rect 162860 79766 162912 79772
rect 163016 79778 163044 80036
rect 163378 79778 163406 80036
rect 163746 79830 163774 80036
rect 160020 75138 160048 75398
rect 160204 75154 160232 79750
rect 160008 75132 160060 75138
rect 160008 75074 160060 75080
rect 160112 75126 160232 75154
rect 160284 75132 160336 75138
rect 158916 64846 159496 64874
rect 158916 49298 158944 64846
rect 158904 49292 158956 49298
rect 158904 49234 158956 49240
rect 160112 27266 160140 75126
rect 160284 75074 160336 75080
rect 160192 75064 160244 75070
rect 160192 75006 160244 75012
rect 160204 50658 160232 75006
rect 160296 64462 160324 75074
rect 160756 75070 160784 79750
rect 160744 75064 160796 75070
rect 160744 75006 160796 75012
rect 160940 65822 160968 79750
rect 160928 65816 160980 65822
rect 160928 65758 160980 65764
rect 160284 64456 160336 64462
rect 160284 64398 160336 64404
rect 160192 50652 160244 50658
rect 160192 50594 160244 50600
rect 160100 27260 160152 27266
rect 160100 27202 160152 27208
rect 161492 27198 161520 79750
rect 161572 75200 161624 75206
rect 161572 75142 161624 75148
rect 161584 28626 161612 75142
rect 161676 52018 161704 79750
rect 162044 67182 162072 79750
rect 162596 75206 162624 79750
rect 162584 75200 162636 75206
rect 162584 75142 162636 75148
rect 162032 67176 162084 67182
rect 162032 67118 162084 67124
rect 161664 52012 161716 52018
rect 161664 51954 161716 51960
rect 162872 41070 162900 79766
rect 163016 79750 163084 79778
rect 162952 75200 163004 75206
rect 162952 75142 163004 75148
rect 162964 53378 162992 75142
rect 163056 53446 163084 79750
rect 163148 79750 163406 79778
rect 163734 79824 163786 79830
rect 164114 79778 164142 80036
rect 163734 79766 163786 79772
rect 164068 79750 164142 79778
rect 164240 79824 164292 79830
rect 164240 79766 164292 79772
rect 164396 79778 164424 80036
rect 164758 79830 164786 80036
rect 164746 79824 164798 79830
rect 163148 68610 163176 79750
rect 164068 75206 164096 79750
rect 164056 75200 164108 75206
rect 164056 75142 164108 75148
rect 163136 68604 163188 68610
rect 163136 68546 163188 68552
rect 163044 53440 163096 53446
rect 163044 53382 163096 53388
rect 162952 53372 163004 53378
rect 162952 53314 163004 53320
rect 162860 41064 162912 41070
rect 162860 41006 162912 41012
rect 161572 28620 161624 28626
rect 161572 28562 161624 28568
rect 164252 28558 164280 79766
rect 164396 79750 164464 79778
rect 165126 79778 165154 80036
rect 164746 79766 164798 79772
rect 164332 75200 164384 75206
rect 164332 75142 164384 75148
rect 164344 54874 164372 75142
rect 164436 69970 164464 79750
rect 165080 79750 165154 79778
rect 165500 79778 165528 80036
rect 165862 79778 165890 80036
rect 166230 79778 166258 80036
rect 165500 79750 165568 79778
rect 165080 75206 165108 79750
rect 165068 75200 165120 75206
rect 165068 75142 165120 75148
rect 165540 71330 165568 79750
rect 165632 79750 165890 79778
rect 166184 79750 166258 79778
rect 166604 79778 166632 80036
rect 166972 79914 167000 80036
rect 166972 79886 167224 79914
rect 167000 79824 167052 79830
rect 166604 79750 166672 79778
rect 167000 79766 167052 79772
rect 165528 71324 165580 71330
rect 165528 71266 165580 71272
rect 164424 69964 164476 69970
rect 164424 69906 164476 69912
rect 164332 54868 164384 54874
rect 164332 54810 164384 54816
rect 165632 29986 165660 79750
rect 166184 70394 166212 79750
rect 166448 78192 166500 78198
rect 166448 78134 166500 78140
rect 165724 70366 166212 70394
rect 165724 56234 165752 70366
rect 166460 64874 166488 78134
rect 166644 72758 166672 79750
rect 166632 72752 166684 72758
rect 166632 72694 166684 72700
rect 166276 64846 166488 64874
rect 165712 56228 165764 56234
rect 165712 56170 165764 56176
rect 165620 29980 165672 29986
rect 165620 29922 165672 29928
rect 164240 28552 164292 28558
rect 164240 28494 164292 28500
rect 161480 27192 161532 27198
rect 161480 27134 161532 27140
rect 160744 27056 160796 27062
rect 160744 26998 160796 27004
rect 158812 22976 158864 22982
rect 158812 22918 158864 22924
rect 160652 14612 160704 14618
rect 160652 14554 160704 14560
rect 158720 13320 158772 13326
rect 158720 13262 158772 13268
rect 157800 13252 157852 13258
rect 157800 13194 157852 13200
rect 155960 11756 156012 11762
rect 155960 11698 156012 11704
rect 156604 3460 156656 3466
rect 156604 3402 156656 3408
rect 156616 480 156644 3402
rect 157812 480 157840 13194
rect 158904 13184 158956 13190
rect 158904 13126 158956 13132
rect 158916 480 158944 13126
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 160664 3482 160692 14554
rect 160756 3670 160784 26998
rect 162124 20120 162176 20126
rect 162124 20062 162176 20068
rect 160836 20052 160888 20058
rect 160836 19994 160888 20000
rect 160744 3664 160796 3670
rect 160744 3606 160796 3612
rect 160848 3602 160876 19994
rect 161480 19984 161532 19990
rect 161480 19926 161532 19932
rect 161492 16574 161520 19926
rect 161492 16546 162072 16574
rect 160836 3596 160888 3602
rect 160836 3538 160888 3544
rect 160112 480 160140 3470
rect 160664 3454 161336 3482
rect 161308 480 161336 3454
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 162136 3738 162164 20062
rect 166276 16114 166304 64846
rect 167012 41002 167040 79766
rect 167196 77382 167224 79886
rect 167334 79778 167362 80036
rect 167702 79778 167730 80036
rect 168070 79830 168098 80036
rect 167288 79750 167362 79778
rect 167472 79750 167730 79778
rect 168058 79824 168110 79830
rect 168058 79766 168110 79772
rect 168444 79778 168472 80036
rect 168812 79778 168840 80036
rect 169174 79778 169202 80036
rect 169542 79778 169570 80036
rect 169758 79928 169814 79937
rect 169916 79914 169944 80036
rect 170278 79937 170306 80036
rect 170264 79928 170320 79937
rect 169916 79886 170076 79914
rect 169758 79863 169814 79872
rect 168444 79750 168604 79778
rect 168812 79750 168880 79778
rect 167184 77376 167236 77382
rect 167184 77318 167236 77324
rect 167288 77194 167316 79750
rect 167104 77166 167316 77194
rect 167104 56166 167132 77166
rect 167472 74118 167500 79750
rect 168472 77308 168524 77314
rect 168472 77250 168524 77256
rect 168380 77240 168432 77246
rect 168380 77182 168432 77188
rect 167460 74112 167512 74118
rect 167460 74054 167512 74060
rect 167092 56160 167144 56166
rect 167092 56102 167144 56108
rect 167000 40996 167052 41002
rect 167000 40938 167052 40944
rect 166356 29776 166408 29782
rect 166356 29718 166408 29724
rect 166264 16108 166316 16114
rect 166264 16050 166316 16056
rect 164424 14544 164476 14550
rect 164424 14486 164476 14492
rect 163688 13116 163740 13122
rect 163688 13058 163740 13064
rect 162124 3732 162176 3738
rect 162124 3674 162176 3680
rect 163700 480 163728 13058
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 14486
rect 166080 6248 166132 6254
rect 166080 6190 166132 6196
rect 166092 480 166120 6190
rect 166368 3466 166396 29718
rect 167000 24200 167052 24206
rect 167000 24142 167052 24148
rect 167012 16574 167040 24142
rect 167012 16546 167224 16574
rect 166356 3460 166408 3466
rect 166356 3402 166408 3408
rect 167196 480 167224 16546
rect 168392 6254 168420 77182
rect 168484 57526 168512 77250
rect 168576 57594 168604 79750
rect 168852 75478 168880 79750
rect 169128 79750 169202 79778
rect 169496 79750 169570 79778
rect 169024 77376 169076 77382
rect 169024 77318 169076 77324
rect 168840 75472 168892 75478
rect 168840 75414 168892 75420
rect 168564 57588 168616 57594
rect 168564 57530 168616 57536
rect 168472 57520 168524 57526
rect 168472 57462 168524 57468
rect 169036 45150 169064 77318
rect 169128 77246 169156 79750
rect 169496 77314 169524 79750
rect 169484 77308 169536 77314
rect 169484 77250 169536 77256
rect 169116 77240 169168 77246
rect 169116 77182 169168 77188
rect 169024 45144 169076 45150
rect 169024 45086 169076 45092
rect 168472 22772 168524 22778
rect 168472 22714 168524 22720
rect 168380 6248 168432 6254
rect 168380 6190 168432 6196
rect 168484 3482 168512 22714
rect 169772 6458 169800 79863
rect 169852 79824 169904 79830
rect 169852 79766 169904 79772
rect 169864 59022 169892 79766
rect 170048 76838 170076 79886
rect 170646 79898 170674 80036
rect 170264 79863 170320 79872
rect 170634 79892 170686 79898
rect 170634 79834 170686 79840
rect 171014 79778 171042 80036
rect 171382 79914 171410 80036
rect 170600 79750 171042 79778
rect 171152 79886 171410 79914
rect 170036 76832 170088 76838
rect 170036 76774 170088 76780
rect 170600 64874 170628 79750
rect 169956 64846 170628 64874
rect 169956 63102 169984 64846
rect 169944 63096 169996 63102
rect 169944 63038 169996 63044
rect 169852 59016 169904 59022
rect 169852 58958 169904 58964
rect 171152 42362 171180 79886
rect 171232 79824 171284 79830
rect 171750 79778 171778 80036
rect 172118 79830 172146 80036
rect 171232 79766 171284 79772
rect 171244 51950 171272 79766
rect 171336 79750 171778 79778
rect 172106 79824 172158 79830
rect 172106 79766 172158 79772
rect 172492 79778 172520 80036
rect 172854 79778 172882 80036
rect 173222 79778 173250 80036
rect 173590 79778 173618 80036
rect 172492 79750 172560 79778
rect 171336 58954 171364 79750
rect 171324 58948 171376 58954
rect 171324 58890 171376 58896
rect 171232 51944 171284 51950
rect 171232 51886 171284 51892
rect 171140 42356 171192 42362
rect 171140 42298 171192 42304
rect 170404 16040 170456 16046
rect 170404 15982 170456 15988
rect 169760 6452 169812 6458
rect 169760 6394 169812 6400
rect 169576 6384 169628 6390
rect 169576 6326 169628 6332
rect 168392 3454 168512 3482
rect 168392 480 168420 3454
rect 169588 480 169616 6326
rect 170416 3806 170444 15982
rect 171968 14476 172020 14482
rect 171968 14418 172020 14424
rect 170404 3800 170456 3806
rect 170404 3742 170456 3748
rect 170772 3596 170824 3602
rect 170772 3538 170824 3544
rect 170784 480 170812 3538
rect 171980 480 172008 14418
rect 172532 6390 172560 79750
rect 172624 79750 172882 79778
rect 172992 79750 173250 79778
rect 173360 79750 173618 79778
rect 173964 79778 173992 80036
rect 174326 79898 174354 80036
rect 174694 79898 174722 80036
rect 174314 79892 174366 79898
rect 174314 79834 174366 79840
rect 174682 79892 174734 79898
rect 174682 79834 174734 79840
rect 175062 79778 175090 80036
rect 175430 79778 175458 80036
rect 175798 79778 175826 80036
rect 176074 79778 176102 80036
rect 176442 79778 176470 80036
rect 173964 79750 174124 79778
rect 172624 13394 172652 79750
rect 172992 77294 173020 79750
rect 172716 77266 173020 77294
rect 172716 20262 172744 77266
rect 173360 64874 173388 79750
rect 173900 79688 173952 79694
rect 173900 79630 173952 79636
rect 173992 79688 174044 79694
rect 173992 79630 174044 79636
rect 172808 64846 173388 64874
rect 172808 29918 172836 64846
rect 172796 29912 172848 29918
rect 172796 29854 172848 29860
rect 172796 21480 172848 21486
rect 172796 21422 172848 21428
rect 172704 20256 172756 20262
rect 172704 20198 172756 20204
rect 172612 13388 172664 13394
rect 172612 13330 172664 13336
rect 172520 6384 172572 6390
rect 172520 6326 172572 6332
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172808 354 172836 21422
rect 173912 20194 173940 79630
rect 174004 31346 174032 79630
rect 174096 60314 174124 79750
rect 174188 79750 175090 79778
rect 175292 79750 175458 79778
rect 175568 79750 175826 79778
rect 176028 79750 176102 79778
rect 176396 79750 176470 79778
rect 176660 79824 176712 79830
rect 176810 79778 176838 80036
rect 177178 79778 177206 80036
rect 177546 79830 177574 80036
rect 176660 79766 176712 79772
rect 174084 60308 174136 60314
rect 174084 60250 174136 60256
rect 174188 60246 174216 79750
rect 174176 60240 174228 60246
rect 174176 60182 174228 60188
rect 173992 31340 174044 31346
rect 173992 31282 174044 31288
rect 174544 31136 174596 31142
rect 174544 31078 174596 31084
rect 173900 20188 173952 20194
rect 173900 20130 173952 20136
rect 174556 3534 174584 31078
rect 175292 20126 175320 79750
rect 175372 77308 175424 77314
rect 175568 77294 175596 79750
rect 175372 77250 175424 77256
rect 175476 77266 175596 77294
rect 175280 20120 175332 20126
rect 175280 20062 175332 20068
rect 175384 20058 175412 77250
rect 175476 31278 175504 77266
rect 176028 64874 176056 79750
rect 176396 77314 176424 79750
rect 176384 77308 176436 77314
rect 176384 77250 176436 77256
rect 175568 64846 176056 64874
rect 175568 60178 175596 64846
rect 175556 60172 175608 60178
rect 175556 60114 175608 60120
rect 175464 31272 175516 31278
rect 175464 31214 175516 31220
rect 175372 20052 175424 20058
rect 175372 19994 175424 20000
rect 175464 15972 175516 15978
rect 175464 15914 175516 15920
rect 174268 3528 174320 3534
rect 174268 3470 174320 3476
rect 174544 3528 174596 3534
rect 174544 3470 174596 3476
rect 174280 480 174308 3470
rect 175476 480 175504 15914
rect 176672 12034 176700 79766
rect 176764 79750 176838 79778
rect 176948 79750 177206 79778
rect 177534 79824 177586 79830
rect 177914 79778 177942 80036
rect 177534 79766 177586 79772
rect 177868 79750 177942 79778
rect 178040 79824 178092 79830
rect 178282 79778 178310 80036
rect 178650 79830 178678 80036
rect 178040 79766 178092 79772
rect 176764 31210 176792 79750
rect 176844 75200 176896 75206
rect 176844 75142 176896 75148
rect 176856 32706 176884 75142
rect 176948 61674 176976 79750
rect 177868 75206 177896 79750
rect 177856 75200 177908 75206
rect 177856 75142 177908 75148
rect 176936 61668 176988 61674
rect 176936 61610 176988 61616
rect 176844 32700 176896 32706
rect 176844 32642 176896 32648
rect 176752 31204 176804 31210
rect 176752 31146 176804 31152
rect 178052 21690 178080 79766
rect 178144 79750 178310 79778
rect 178638 79824 178690 79830
rect 179018 79778 179046 80036
rect 178638 79766 178690 79772
rect 178788 79750 179046 79778
rect 179392 79778 179420 80036
rect 179754 79778 179782 80036
rect 180122 79778 180150 80036
rect 180490 79778 180518 80036
rect 179392 79750 179460 79778
rect 178144 61606 178172 79750
rect 178788 64874 178816 79750
rect 179432 75426 179460 79750
rect 179340 75398 179460 75426
rect 179524 79750 179782 79778
rect 180076 79750 180150 79778
rect 180260 79750 180518 79778
rect 180864 79778 180892 80036
rect 181226 79778 181254 80036
rect 181594 79778 181622 80036
rect 181962 79778 181990 80036
rect 180864 79750 180932 79778
rect 179340 75138 179368 75398
rect 179524 75154 179552 79750
rect 179328 75132 179380 75138
rect 179328 75074 179380 75080
rect 179432 75126 179552 75154
rect 179604 75132 179656 75138
rect 178236 64846 178816 64874
rect 178132 61600 178184 61606
rect 178132 61542 178184 61548
rect 178132 50380 178184 50386
rect 178132 50322 178184 50328
rect 178040 21684 178092 21690
rect 178040 21626 178092 21632
rect 176752 21412 176804 21418
rect 176752 21354 176804 21360
rect 176660 12028 176712 12034
rect 176660 11970 176712 11976
rect 176764 6914 176792 21354
rect 178144 16574 178172 50322
rect 178236 32638 178264 64846
rect 178224 32632 178276 32638
rect 178224 32574 178276 32580
rect 179432 18902 179460 75126
rect 179604 75074 179656 75080
rect 179512 75064 179564 75070
rect 179512 75006 179564 75012
rect 179524 32570 179552 75006
rect 179616 61538 179644 75074
rect 180076 75070 180104 79750
rect 180064 75064 180116 75070
rect 180064 75006 180116 75012
rect 180260 64874 180288 79750
rect 180800 75200 180852 75206
rect 180800 75142 180852 75148
rect 179708 64846 180288 64874
rect 179708 63034 179736 64846
rect 179696 63028 179748 63034
rect 179696 62970 179748 62976
rect 179604 61532 179656 61538
rect 179604 61474 179656 61480
rect 179512 32564 179564 32570
rect 179512 32506 179564 32512
rect 179512 21548 179564 21554
rect 179512 21490 179564 21496
rect 179420 18896 179472 18902
rect 179420 18838 179472 18844
rect 179524 16574 179552 21490
rect 178144 16546 178632 16574
rect 179524 16546 180288 16574
rect 176672 6886 176792 6914
rect 176672 480 176700 6886
rect 177856 3596 177908 3602
rect 177856 3538 177908 3544
rect 177868 480 177896 3538
rect 173134 354 173246 480
rect 172808 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 180812 5098 180840 75142
rect 180904 17542 180932 79750
rect 180996 79750 181254 79778
rect 181548 79750 181622 79778
rect 181916 79750 181990 79778
rect 182180 79824 182232 79830
rect 182330 79778 182358 80036
rect 182698 79778 182726 80036
rect 183066 79830 183094 80036
rect 182180 79766 182232 79772
rect 180996 34066 181024 79750
rect 181548 64874 181576 79750
rect 181916 75206 181944 79750
rect 181904 75200 181956 75206
rect 181904 75142 181956 75148
rect 181088 64846 181576 64874
rect 181088 62966 181116 64846
rect 181076 62960 181128 62966
rect 181076 62902 181128 62908
rect 181076 40792 181128 40798
rect 181076 40734 181128 40740
rect 180984 34060 181036 34066
rect 180984 34002 181036 34008
rect 180892 17536 180944 17542
rect 180892 17478 180944 17484
rect 180800 5092 180852 5098
rect 180800 5034 180852 5040
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181088 354 181116 40734
rect 182192 21622 182220 79766
rect 182284 79750 182358 79778
rect 182468 79750 182726 79778
rect 183054 79824 183106 79830
rect 183434 79778 183462 80036
rect 183652 79892 183704 79898
rect 183652 79834 183704 79840
rect 183054 79766 183106 79772
rect 183388 79750 183462 79778
rect 183560 79824 183612 79830
rect 183560 79766 183612 79772
rect 182284 33998 182312 79750
rect 182364 75200 182416 75206
rect 182364 75142 182416 75148
rect 182272 33992 182324 33998
rect 182272 33934 182324 33940
rect 182376 33930 182404 75142
rect 182468 62898 182496 79750
rect 183388 75206 183416 79750
rect 183376 75200 183428 75206
rect 183376 75142 183428 75148
rect 182456 62892 182508 62898
rect 182456 62834 182508 62840
rect 182364 33924 182416 33930
rect 182364 33866 182416 33872
rect 182180 21616 182232 21622
rect 182180 21558 182232 21564
rect 183572 21554 183600 79766
rect 183664 35426 183692 79834
rect 183802 79778 183830 80036
rect 184170 79830 184198 80036
rect 184538 79898 184566 80036
rect 184526 79892 184578 79898
rect 184526 79834 184578 79840
rect 183756 79750 183830 79778
rect 184158 79824 184210 79830
rect 184158 79766 184210 79772
rect 184912 79778 184940 80036
rect 185274 79778 185302 80036
rect 184912 79750 184980 79778
rect 183756 64394 183784 79750
rect 184952 75426 184980 79750
rect 184860 75398 184980 75426
rect 185044 79750 185302 79778
rect 185648 79778 185676 80036
rect 186010 79778 186038 80036
rect 186378 79778 186406 80036
rect 186746 79778 186774 80036
rect 187114 79778 187142 80036
rect 185648 79750 185716 79778
rect 184860 75138 184888 75398
rect 185044 75154 185072 79750
rect 185688 78538 185716 79750
rect 185964 79750 186038 79778
rect 186332 79750 186406 79778
rect 186516 79750 186774 79778
rect 186884 79750 187142 79778
rect 187488 79778 187516 80036
rect 187850 79914 187878 80036
rect 187712 79886 187878 79914
rect 187488 79750 187556 79778
rect 185676 78532 185728 78538
rect 185676 78474 185728 78480
rect 184848 75132 184900 75138
rect 184848 75074 184900 75080
rect 184952 75126 185072 75154
rect 185124 75132 185176 75138
rect 183744 64388 183796 64394
rect 183744 64330 183796 64336
rect 184204 44940 184256 44946
rect 184204 44882 184256 44888
rect 183652 35420 183704 35426
rect 183652 35362 183704 35368
rect 183652 24132 183704 24138
rect 183652 24074 183704 24080
rect 183560 21548 183612 21554
rect 183560 21490 183612 21496
rect 183664 16574 183692 24074
rect 183664 16546 183784 16574
rect 182180 16108 182232 16114
rect 182180 16050 182232 16056
rect 181414 354 181526 480
rect 181088 326 181526 354
rect 182192 354 182220 16050
rect 183756 480 183784 16546
rect 184216 2990 184244 44882
rect 184952 21486 184980 75126
rect 185124 75074 185176 75080
rect 185032 75064 185084 75070
rect 185032 75006 185084 75012
rect 185044 64258 185072 75006
rect 185136 64326 185164 75074
rect 185964 75070 185992 79750
rect 185952 75064 186004 75070
rect 185952 75006 186004 75012
rect 185124 64320 185176 64326
rect 185124 64262 185176 64268
rect 185032 64252 185084 64258
rect 185032 64194 185084 64200
rect 185032 28348 185084 28354
rect 185032 28290 185084 28296
rect 184940 21480 184992 21486
rect 184940 21422 184992 21428
rect 185044 6914 185072 28290
rect 186332 25770 186360 79750
rect 186516 77330 186544 79750
rect 186424 77302 186544 77330
rect 186424 36854 186452 77302
rect 186884 65754 186912 79750
rect 187056 78056 187108 78062
rect 187056 77998 187108 78004
rect 186964 77988 187016 77994
rect 186964 77930 187016 77936
rect 186872 65748 186924 65754
rect 186872 65690 186924 65696
rect 186412 36848 186464 36854
rect 186412 36790 186464 36796
rect 186320 25764 186372 25770
rect 186320 25706 186372 25712
rect 184952 6886 185072 6914
rect 184204 2984 184256 2990
rect 184204 2926 184256 2932
rect 184952 480 184980 6886
rect 186136 3664 186188 3670
rect 186136 3606 186188 3612
rect 186148 480 186176 3606
rect 186976 3602 187004 77930
rect 187068 5166 187096 77998
rect 187528 77450 187556 79750
rect 187516 77444 187568 77450
rect 187516 77386 187568 77392
rect 187712 7886 187740 79886
rect 187792 79824 187844 79830
rect 188126 79778 188154 80036
rect 187792 79766 187844 79772
rect 187700 7880 187752 7886
rect 187700 7822 187752 7828
rect 187804 7818 187832 79766
rect 187896 79750 188154 79778
rect 188500 79778 188528 80036
rect 188862 79830 188890 80036
rect 189080 79892 189132 79898
rect 189080 79834 189132 79840
rect 188850 79824 188902 79830
rect 188500 79750 188568 79778
rect 188850 79766 188902 79772
rect 187896 65686 187924 79750
rect 188540 78606 188568 79750
rect 188528 78600 188580 78606
rect 188528 78542 188580 78548
rect 188344 78124 188396 78130
rect 188344 78066 188396 78072
rect 187884 65680 187936 65686
rect 187884 65622 187936 65628
rect 188356 18834 188384 78066
rect 189092 45082 189120 79834
rect 189230 79778 189258 80036
rect 189184 79750 189258 79778
rect 189604 79778 189632 80036
rect 189966 79898 189994 80036
rect 189954 79892 190006 79898
rect 189954 79834 190006 79840
rect 190334 79778 190362 80036
rect 190708 79914 190736 80036
rect 190708 79886 190776 79914
rect 189604 79750 189672 79778
rect 189184 65618 189212 79750
rect 189644 78674 189672 79750
rect 189736 79750 190362 79778
rect 190460 79824 190512 79830
rect 190460 79766 190512 79772
rect 189632 78668 189684 78674
rect 189632 78610 189684 78616
rect 189736 67114 189764 79750
rect 189724 67108 189776 67114
rect 189724 67050 189776 67056
rect 189172 65612 189224 65618
rect 189172 65554 189224 65560
rect 189080 45076 189132 45082
rect 189080 45018 189132 45024
rect 188436 35352 188488 35358
rect 188436 35294 188488 35300
rect 188344 18828 188396 18834
rect 188344 18770 188396 18776
rect 187792 7812 187844 7818
rect 187792 7754 187844 7760
rect 187332 7676 187384 7682
rect 187332 7618 187384 7624
rect 187056 5160 187108 5166
rect 187056 5102 187108 5108
rect 186964 3596 187016 3602
rect 186964 3538 187016 3544
rect 187344 480 187372 7618
rect 188448 3738 188476 35294
rect 190472 7750 190500 79766
rect 190748 77722 190776 79886
rect 191070 79830 191098 80036
rect 191058 79824 191110 79830
rect 191438 79778 191466 80036
rect 191058 79766 191110 79772
rect 191208 79750 191466 79778
rect 191812 79778 191840 80036
rect 192174 79778 192202 80036
rect 192542 79778 192570 80036
rect 191812 79750 191880 79778
rect 190736 77716 190788 77722
rect 190736 77658 190788 77664
rect 191208 77602 191236 79750
rect 191380 78668 191432 78674
rect 191380 78610 191432 78616
rect 191288 78532 191340 78538
rect 191288 78474 191340 78480
rect 190564 77574 191236 77602
rect 190564 14754 190592 77574
rect 191300 77466 191328 78474
rect 191104 77444 191156 77450
rect 191104 77386 191156 77392
rect 191208 77438 191328 77466
rect 190644 25560 190696 25566
rect 190644 25502 190696 25508
rect 190552 14748 190604 14754
rect 190552 14690 190604 14696
rect 188528 7744 188580 7750
rect 188528 7686 188580 7692
rect 190460 7744 190512 7750
rect 190460 7686 190512 7692
rect 188436 3732 188488 3738
rect 188436 3674 188488 3680
rect 188540 480 188568 7686
rect 189724 2984 189776 2990
rect 189724 2926 189776 2932
rect 189736 480 189764 2926
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190656 354 190684 25502
rect 191116 16182 191144 77386
rect 191208 35494 191236 77438
rect 191392 64874 191420 78610
rect 191852 77314 191880 79750
rect 191944 79750 192202 79778
rect 192496 79750 192570 79778
rect 192916 79778 192944 80036
rect 193284 79778 193312 80036
rect 193404 79824 193456 79830
rect 192916 79750 192984 79778
rect 193284 79750 193352 79778
rect 193646 79778 193674 80036
rect 194020 79914 194048 80036
rect 194020 79886 194088 79914
rect 193404 79766 193456 79772
rect 191840 77308 191892 77314
rect 191840 77250 191892 77256
rect 191840 77172 191892 77178
rect 191840 77114 191892 77120
rect 191300 64846 191420 64874
rect 191300 49230 191328 64846
rect 191288 49224 191340 49230
rect 191288 49166 191340 49172
rect 191196 35488 191248 35494
rect 191196 35430 191248 35436
rect 191104 16176 191156 16182
rect 191104 16118 191156 16124
rect 191852 14686 191880 77114
rect 191944 36786 191972 79750
rect 192392 77716 192444 77722
rect 192392 77658 192444 77664
rect 192024 77308 192076 77314
rect 192024 77250 192076 77256
rect 192036 46442 192064 77250
rect 192404 74534 192432 77658
rect 192496 77178 192524 79750
rect 192576 78600 192628 78606
rect 192576 78542 192628 78548
rect 192484 77172 192536 77178
rect 192484 77114 192536 77120
rect 192404 74506 192524 74534
rect 192024 46436 192076 46442
rect 192024 46378 192076 46384
rect 191932 36780 191984 36786
rect 191932 36722 191984 36728
rect 191840 14680 191892 14686
rect 191840 14622 191892 14628
rect 192496 10606 192524 74506
rect 192588 28490 192616 78542
rect 192956 77382 192984 79750
rect 192944 77376 192996 77382
rect 192944 77318 192996 77324
rect 193220 77308 193272 77314
rect 193220 77250 193272 77256
rect 192576 28484 192628 28490
rect 192576 28426 192628 28432
rect 193232 14618 193260 77250
rect 193324 36718 193352 79750
rect 193416 45014 193444 79766
rect 193600 79750 193674 79778
rect 193600 77314 193628 79750
rect 194060 77382 194088 79886
rect 194382 79830 194410 80036
rect 194370 79824 194422 79830
rect 194370 79766 194422 79772
rect 194600 79824 194652 79830
rect 194600 79766 194652 79772
rect 194756 79778 194784 80036
rect 195118 79778 195146 80036
rect 195486 79830 195514 80036
rect 193864 77376 193916 77382
rect 193864 77318 193916 77324
rect 194048 77376 194100 77382
rect 194048 77318 194100 77324
rect 193588 77308 193640 77314
rect 193588 77250 193640 77256
rect 193404 45008 193456 45014
rect 193404 44950 193456 44956
rect 193876 42294 193904 77318
rect 193864 42288 193916 42294
rect 193864 42230 193916 42236
rect 194612 38214 194640 79766
rect 194756 79750 194824 79778
rect 194692 77308 194744 77314
rect 194692 77250 194744 77256
rect 194704 61470 194732 77250
rect 194796 67046 194824 79750
rect 195072 79750 195146 79778
rect 195474 79824 195526 79830
rect 195474 79766 195526 79772
rect 195860 79778 195888 80036
rect 196222 79778 196250 80036
rect 196590 79778 196618 80036
rect 196958 79778 196986 80036
rect 195860 79750 195928 79778
rect 195072 77314 195100 79750
rect 195244 77376 195296 77382
rect 195244 77318 195296 77324
rect 195060 77308 195112 77314
rect 195060 77250 195112 77256
rect 194784 67040 194836 67046
rect 194784 66982 194836 66988
rect 194692 61464 194744 61470
rect 194692 61406 194744 61412
rect 195256 50590 195284 77318
rect 195900 75410 195928 79750
rect 195992 79750 196250 79778
rect 196360 79750 196618 79778
rect 196728 79750 196986 79778
rect 197332 79778 197360 80036
rect 197694 79778 197722 80036
rect 198062 79778 198090 80036
rect 197332 79750 197400 79778
rect 195888 75404 195940 75410
rect 195888 75346 195940 75352
rect 195244 50584 195296 50590
rect 195244 50526 195296 50532
rect 194600 38208 194652 38214
rect 194600 38150 194652 38156
rect 193312 36712 193364 36718
rect 193312 36654 193364 36660
rect 195992 29850 196020 79750
rect 196360 77330 196388 79750
rect 196084 77302 196388 77330
rect 196084 46374 196112 77302
rect 196728 72690 196756 79750
rect 196716 72684 196768 72690
rect 196716 72626 196768 72632
rect 196072 46368 196124 46374
rect 196072 46310 196124 46316
rect 195980 29844 196032 29850
rect 195980 29786 196032 29792
rect 197372 27130 197400 79750
rect 197464 79750 197722 79778
rect 197832 79750 198090 79778
rect 198436 79778 198464 80036
rect 198804 79778 198832 80036
rect 198924 79824 198976 79830
rect 198436 79750 198504 79778
rect 198804 79750 198872 79778
rect 199166 79778 199194 80036
rect 199534 79778 199562 80036
rect 199902 79830 199930 80036
rect 198924 79766 198976 79772
rect 197464 38146 197492 79750
rect 197832 69902 197860 79750
rect 198476 78062 198504 79750
rect 198464 78056 198516 78062
rect 198464 77998 198516 78004
rect 198740 77308 198792 77314
rect 198740 77250 198792 77256
rect 197820 69896 197872 69902
rect 197820 69838 197872 69844
rect 197452 38140 197504 38146
rect 197452 38082 197504 38088
rect 197452 28280 197504 28286
rect 197452 28222 197504 28228
rect 197360 27124 197412 27130
rect 197360 27066 197412 27072
rect 193312 26988 193364 26994
rect 193312 26930 193364 26936
rect 193220 14612 193272 14618
rect 193220 14554 193272 14560
rect 192484 10600 192536 10606
rect 192484 10542 192536 10548
rect 193324 3670 193352 26930
rect 195980 17400 196032 17406
rect 195980 17342 196032 17348
rect 195992 16574 196020 17342
rect 197464 16574 197492 28222
rect 195992 16546 196848 16574
rect 197464 16546 197952 16574
rect 193404 15904 193456 15910
rect 193404 15846 193456 15852
rect 193312 3664 193364 3670
rect 193312 3606 193364 3612
rect 193416 3482 193444 15846
rect 194416 3664 194468 3670
rect 194416 3606 194468 3612
rect 192024 3460 192076 3466
rect 192024 3402 192076 3408
rect 193232 3454 193444 3482
rect 192036 480 192064 3402
rect 193232 480 193260 3454
rect 194428 480 194456 3606
rect 195612 3528 195664 3534
rect 195612 3470 195664 3476
rect 195624 480 195652 3470
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 198752 9246 198780 77250
rect 198844 38078 198872 79750
rect 198936 39642 198964 79766
rect 199028 79750 199194 79778
rect 199488 79750 199562 79778
rect 199890 79824 199942 79830
rect 199890 79766 199942 79772
rect 200184 79778 200212 80036
rect 200546 79898 200574 80036
rect 200914 79898 200942 80036
rect 200534 79892 200586 79898
rect 200534 79834 200586 79840
rect 200902 79892 200954 79898
rect 200902 79834 200954 79840
rect 201282 79778 201310 80036
rect 201656 79914 201684 80036
rect 201656 79886 201724 79914
rect 200184 79750 200344 79778
rect 199028 68542 199056 79750
rect 199488 77314 199516 79750
rect 200120 79688 200172 79694
rect 200120 79630 200172 79636
rect 200212 79688 200264 79694
rect 200212 79630 200264 79636
rect 199476 77308 199528 77314
rect 199476 77250 199528 77256
rect 199016 68536 199068 68542
rect 199016 68478 199068 68484
rect 198924 39636 198976 39642
rect 198924 39578 198976 39584
rect 198832 38072 198884 38078
rect 198832 38014 198884 38020
rect 200132 14550 200160 79630
rect 200224 39574 200252 79630
rect 200316 66978 200344 79750
rect 200408 79750 201310 79778
rect 200408 68474 200436 79750
rect 201696 77518 201724 79886
rect 202018 79778 202046 80036
rect 202386 79778 202414 80036
rect 201788 79750 202046 79778
rect 202156 79750 202414 79778
rect 202760 79778 202788 80036
rect 203122 79778 203150 80036
rect 203490 79778 203518 80036
rect 202760 79750 202828 79778
rect 201684 77512 201736 77518
rect 201684 77454 201736 77460
rect 201788 77330 201816 79750
rect 201512 77302 201816 77330
rect 200396 68468 200448 68474
rect 200396 68410 200448 68416
rect 200304 66972 200356 66978
rect 200304 66914 200356 66920
rect 200212 39568 200264 39574
rect 200212 39510 200264 39516
rect 200212 17332 200264 17338
rect 200212 17274 200264 17280
rect 200224 16574 200252 17274
rect 200224 16546 200344 16574
rect 200120 14544 200172 14550
rect 200120 14486 200172 14492
rect 198740 9240 198792 9246
rect 198740 9182 198792 9188
rect 199108 3732 199160 3738
rect 199108 3674 199160 3680
rect 199120 480 199148 3674
rect 200316 480 200344 16546
rect 201512 9178 201540 77302
rect 202156 68406 202184 79750
rect 202800 77450 202828 79750
rect 202892 79750 203150 79778
rect 203444 79750 203518 79778
rect 203864 79778 203892 80036
rect 204232 79778 204260 80036
rect 204352 79824 204404 79830
rect 203864 79750 203932 79778
rect 204232 79750 204300 79778
rect 204594 79778 204622 80036
rect 204352 79766 204404 79772
rect 202788 77444 202840 77450
rect 202788 77386 202840 77392
rect 202144 68400 202196 68406
rect 202144 68342 202196 68348
rect 202892 40934 202920 79750
rect 203444 69834 203472 79750
rect 203524 78056 203576 78062
rect 203524 77998 203576 78004
rect 203432 69828 203484 69834
rect 203432 69770 203484 69776
rect 202880 40928 202932 40934
rect 202880 40870 202932 40876
rect 201592 29708 201644 29714
rect 201592 29650 201644 29656
rect 201500 9172 201552 9178
rect 201500 9114 201552 9120
rect 201604 6914 201632 29650
rect 202880 17264 202932 17270
rect 202880 17206 202932 17212
rect 202892 16574 202920 17206
rect 202892 16546 203472 16574
rect 202696 9036 202748 9042
rect 202696 8978 202748 8984
rect 201512 6886 201632 6914
rect 201512 480 201540 6886
rect 202708 480 202736 8978
rect 190798 354 190910 480
rect 190656 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 203536 6322 203564 77998
rect 203904 77314 203932 79750
rect 203892 77308 203944 77314
rect 203892 77250 203944 77256
rect 204272 39438 204300 79750
rect 204364 46306 204392 79766
rect 204456 79750 204622 79778
rect 204968 79778 204996 80036
rect 205330 79830 205358 80036
rect 205318 79824 205370 79830
rect 204968 79750 205036 79778
rect 205318 79766 205370 79772
rect 205704 79778 205732 80036
rect 206072 79914 206100 80036
rect 206072 79886 206140 79914
rect 206434 79898 206462 80036
rect 205704 79750 205772 79778
rect 204456 69766 204484 79750
rect 205008 78538 205036 79750
rect 205640 79688 205692 79694
rect 205640 79630 205692 79636
rect 204996 78532 205048 78538
rect 204996 78474 205048 78480
rect 204444 69760 204496 69766
rect 204444 69702 204496 69708
rect 204352 46300 204404 46306
rect 204352 46242 204404 46248
rect 204260 39432 204312 39438
rect 204260 39374 204312 39380
rect 204260 29640 204312 29646
rect 204260 29582 204312 29588
rect 204272 16574 204300 29582
rect 204272 16546 205128 16574
rect 203524 6316 203576 6322
rect 203524 6258 203576 6264
rect 205100 480 205128 16546
rect 205652 9110 205680 79630
rect 205744 16114 205772 79750
rect 206112 77382 206140 79886
rect 206422 79892 206474 79898
rect 206422 79834 206474 79840
rect 206802 79778 206830 80036
rect 207176 79914 207204 80036
rect 207176 79886 207244 79914
rect 206204 79750 206830 79778
rect 206100 77376 206152 77382
rect 206100 77318 206152 77324
rect 206204 64874 206232 79750
rect 207216 78266 207244 79886
rect 207538 79778 207566 80036
rect 207906 79778 207934 80036
rect 207308 79750 207566 79778
rect 207676 79750 207934 79778
rect 208280 79778 208308 80036
rect 208400 79824 208452 79830
rect 208280 79750 208348 79778
rect 208642 79778 208670 80036
rect 209010 79830 209038 80036
rect 208400 79766 208452 79772
rect 207204 78260 207256 78266
rect 207204 78202 207256 78208
rect 207308 77466 207336 79750
rect 207032 77438 207336 77466
rect 206284 77308 206336 77314
rect 206284 77250 206336 77256
rect 205836 64846 206232 64874
rect 205732 16108 205784 16114
rect 205732 16050 205784 16056
rect 205836 16046 205864 64846
rect 206296 39506 206324 77250
rect 207032 46238 207060 77438
rect 207676 77330 207704 79750
rect 208320 78062 208348 79750
rect 208308 78056 208360 78062
rect 208308 77998 208360 78004
rect 207756 77444 207808 77450
rect 207756 77386 207808 77392
rect 207124 77302 207704 77330
rect 207124 71262 207152 77302
rect 207112 71256 207164 71262
rect 207112 71198 207164 71204
rect 207768 64874 207796 77386
rect 207676 64846 207796 64874
rect 207020 46232 207072 46238
rect 207020 46174 207072 46180
rect 206284 39500 206336 39506
rect 206284 39442 206336 39448
rect 207676 19990 207704 64846
rect 207664 19984 207716 19990
rect 207664 19926 207716 19932
rect 205824 16040 205876 16046
rect 205824 15982 205876 15988
rect 208412 15978 208440 79766
rect 208504 79750 208670 79778
rect 208998 79824 209050 79830
rect 208998 79766 209050 79772
rect 209384 79778 209412 80036
rect 209752 79914 209780 80036
rect 209752 79886 209912 79914
rect 209780 79824 209832 79830
rect 209384 79750 209452 79778
rect 209780 79766 209832 79772
rect 208504 42226 208532 79750
rect 209424 78130 209452 79750
rect 209412 78124 209464 78130
rect 209412 78066 209464 78072
rect 209044 77512 209096 77518
rect 209044 77454 209096 77460
rect 208492 42220 208544 42226
rect 208492 42162 208544 42168
rect 208492 31068 208544 31074
rect 208492 31010 208544 31016
rect 208504 16574 208532 31010
rect 208504 16546 208624 16574
rect 208400 15972 208452 15978
rect 208400 15914 208452 15920
rect 205640 9104 205692 9110
rect 205640 9046 205692 9052
rect 206192 8968 206244 8974
rect 206192 8910 206244 8916
rect 206204 480 206232 8910
rect 207388 3596 207440 3602
rect 207388 3538 207440 3544
rect 207400 480 207428 3538
rect 208596 480 208624 16546
rect 209056 7682 209084 77454
rect 209136 77376 209188 77382
rect 209136 77318 209188 77324
rect 209148 31142 209176 77318
rect 209136 31136 209188 31142
rect 209136 31078 209188 31084
rect 209792 12866 209820 79766
rect 209884 42158 209912 79886
rect 210114 79778 210142 80036
rect 209976 79750 210142 79778
rect 210488 79778 210516 80036
rect 210850 79830 210878 80036
rect 210838 79824 210890 79830
rect 210488 79750 210556 79778
rect 210838 79766 210890 79772
rect 211224 79778 211252 80036
rect 211586 79778 211614 80036
rect 211954 79914 211982 80036
rect 211224 79750 211384 79778
rect 209976 71194 210004 79750
rect 210424 78532 210476 78538
rect 210424 78474 210476 78480
rect 209964 71188 210016 71194
rect 209964 71130 210016 71136
rect 209872 42152 209924 42158
rect 209872 42094 209924 42100
rect 209872 40724 209924 40730
rect 209872 40666 209924 40672
rect 209884 16574 209912 40666
rect 210436 21418 210464 78474
rect 210528 77382 210556 79750
rect 210516 77376 210568 77382
rect 210516 77318 210568 77324
rect 211252 77308 211304 77314
rect 211252 77250 211304 77256
rect 211160 77240 211212 77246
rect 211160 77182 211212 77188
rect 210516 44872 210568 44878
rect 210516 44814 210568 44820
rect 210424 21412 210476 21418
rect 210424 21354 210476 21360
rect 209884 16546 210464 16574
rect 209792 12838 209912 12866
rect 209780 9308 209832 9314
rect 209780 9250 209832 9256
rect 209044 7676 209096 7682
rect 209044 7618 209096 7624
rect 209792 480 209820 9250
rect 209884 9042 209912 12838
rect 209872 9036 209924 9042
rect 209872 8978 209924 8984
rect 210436 3482 210464 16546
rect 210528 3602 210556 44814
rect 211172 43722 211200 77182
rect 211264 44946 211292 77250
rect 211356 71126 211384 79750
rect 211540 79750 211614 79778
rect 211724 79886 211982 79914
rect 211540 77314 211568 79750
rect 211528 77308 211580 77314
rect 211528 77250 211580 77256
rect 211724 77246 211752 79886
rect 212230 79778 212258 80036
rect 212598 79778 212626 80036
rect 212966 79778 212994 80036
rect 213334 79778 213362 80036
rect 211816 79750 212258 79778
rect 212552 79750 212626 79778
rect 212736 79750 212994 79778
rect 213288 79750 213362 79778
rect 213708 79778 213736 80036
rect 213920 79824 213972 79830
rect 213708 79750 213776 79778
rect 214070 79778 214098 80036
rect 214444 79914 214472 80036
rect 214444 79886 214512 79914
rect 213920 79766 213972 79772
rect 211712 77240 211764 77246
rect 211712 77182 211764 77188
rect 211816 72622 211844 79750
rect 211804 72616 211856 72622
rect 211804 72558 211856 72564
rect 211344 71120 211396 71126
rect 211344 71062 211396 71068
rect 211252 44940 211304 44946
rect 211252 44882 211304 44888
rect 211160 43716 211212 43722
rect 211160 43658 211212 43664
rect 212552 24410 212580 79750
rect 212632 77308 212684 77314
rect 212632 77250 212684 77256
rect 212644 74050 212672 77250
rect 212632 74044 212684 74050
rect 212632 73986 212684 73992
rect 212736 43586 212764 79750
rect 213092 78260 213144 78266
rect 213092 78202 213144 78208
rect 213104 74534 213132 78202
rect 213184 78056 213236 78062
rect 213184 77998 213236 78004
rect 213196 77194 213224 77998
rect 213288 77314 213316 79750
rect 213748 77314 213776 79750
rect 213276 77308 213328 77314
rect 213276 77250 213328 77256
rect 213736 77308 213788 77314
rect 213736 77250 213788 77256
rect 213196 77166 213316 77194
rect 213104 74506 213224 74534
rect 212724 43580 212776 43586
rect 212724 43522 212776 43528
rect 212632 43444 212684 43450
rect 212632 43386 212684 43392
rect 212540 24404 212592 24410
rect 212540 24346 212592 24352
rect 212644 16574 212672 43386
rect 213196 32502 213224 74506
rect 213288 33862 213316 77166
rect 213276 33856 213328 33862
rect 213276 33798 213328 33804
rect 213184 32496 213236 32502
rect 213184 32438 213236 32444
rect 212644 16546 213408 16574
rect 210516 3596 210568 3602
rect 210516 3538 210568 3544
rect 212172 3596 212224 3602
rect 212172 3538 212224 3544
rect 210436 3454 211016 3482
rect 210988 480 211016 3454
rect 212184 480 212212 3538
rect 213380 480 213408 16546
rect 213932 5030 213960 79766
rect 214024 79750 214098 79778
rect 214024 43518 214052 79750
rect 214104 77240 214156 77246
rect 214104 77182 214156 77188
rect 214116 53310 214144 77182
rect 214484 75342 214512 79886
rect 214806 79778 214834 80036
rect 215174 79830 215202 80036
rect 215548 79914 215576 80036
rect 215916 79914 215944 80036
rect 215548 79886 215616 79914
rect 215916 79886 215984 79914
rect 214760 79750 214834 79778
rect 215162 79824 215214 79830
rect 215162 79766 215214 79772
rect 214564 78124 214616 78130
rect 214564 78066 214616 78072
rect 214472 75336 214524 75342
rect 214472 75278 214524 75284
rect 214104 53304 214156 53310
rect 214104 53246 214156 53252
rect 214012 43512 214064 43518
rect 214012 43454 214064 43460
rect 214576 36650 214604 78066
rect 214760 77246 214788 79750
rect 214748 77240 214800 77246
rect 214748 77182 214800 77188
rect 215588 75274 215616 79886
rect 215956 78198 215984 79886
rect 216278 79778 216306 80036
rect 216652 79914 216680 80036
rect 216652 79886 216812 79914
rect 216048 79750 216306 79778
rect 215944 78192 215996 78198
rect 215944 78134 215996 78140
rect 216048 77466 216076 79750
rect 215772 77438 216076 77466
rect 215576 75268 215628 75274
rect 215576 75210 215628 75216
rect 215772 64874 215800 77438
rect 215944 77308 215996 77314
rect 215944 77250 215996 77256
rect 215312 64846 215800 64874
rect 215312 47802 215340 64846
rect 215300 47796 215352 47802
rect 215300 47738 215352 47744
rect 215956 43654 215984 77250
rect 216784 76770 216812 79886
rect 217014 79778 217042 80036
rect 217382 79778 217410 80036
rect 216876 79750 217042 79778
rect 217244 79750 217410 79778
rect 217756 79778 217784 80036
rect 218124 79778 218152 80036
rect 218486 79778 218514 80036
rect 218854 79778 218882 80036
rect 219222 79778 219250 80036
rect 217756 79750 217824 79778
rect 218124 79750 218192 79778
rect 216772 76764 216824 76770
rect 216772 76706 216824 76712
rect 216876 76650 216904 79750
rect 216692 76622 216904 76650
rect 215944 43648 215996 43654
rect 215944 43590 215996 43596
rect 216692 40866 216720 76622
rect 217244 64874 217272 79750
rect 217324 77376 217376 77382
rect 217324 77318 217376 77324
rect 216784 64846 217272 64874
rect 216784 47734 216812 64846
rect 216772 47728 216824 47734
rect 216772 47670 216824 47676
rect 216680 40860 216732 40866
rect 216680 40802 216732 40808
rect 217336 38010 217364 77318
rect 217796 76702 217824 79750
rect 218164 77314 218192 79750
rect 218256 79750 218514 79778
rect 218808 79750 218882 79778
rect 219176 79750 219250 79778
rect 219440 79824 219492 79830
rect 219440 79766 219492 79772
rect 219596 79778 219624 80036
rect 219958 79830 219986 80036
rect 219946 79824 219998 79830
rect 218152 77308 218204 77314
rect 218152 77250 218204 77256
rect 218060 77240 218112 77246
rect 218060 77182 218112 77188
rect 217784 76696 217836 76702
rect 217784 76638 217836 76644
rect 217324 38004 217376 38010
rect 217324 37946 217376 37952
rect 214564 36644 214616 36650
rect 214564 36586 214616 36592
rect 215300 32428 215352 32434
rect 215300 32370 215352 32376
rect 214012 18760 214064 18766
rect 214012 18702 214064 18708
rect 214024 16574 214052 18702
rect 214024 16546 214512 16574
rect 213920 5024 213972 5030
rect 213920 4966 213972 4972
rect 214484 480 214512 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 32370
rect 218072 22914 218100 77182
rect 218152 77172 218204 77178
rect 218152 77114 218204 77120
rect 218164 32434 218192 77114
rect 218256 47666 218284 79750
rect 218336 77308 218388 77314
rect 218336 77250 218388 77256
rect 218348 54806 218376 77250
rect 218808 77178 218836 79750
rect 219176 77246 219204 79750
rect 219164 77240 219216 77246
rect 219164 77182 219216 77188
rect 218796 77172 218848 77178
rect 218796 77114 218848 77120
rect 218336 54800 218388 54806
rect 218336 54742 218388 54748
rect 218244 47660 218296 47666
rect 218244 47602 218296 47608
rect 218244 33788 218296 33794
rect 218244 33730 218296 33736
rect 218152 32428 218204 32434
rect 218152 32370 218204 32376
rect 218060 22908 218112 22914
rect 218060 22850 218112 22856
rect 218256 16574 218284 33730
rect 218256 16546 219296 16574
rect 216864 10396 216916 10402
rect 216864 10338 216916 10344
rect 216876 480 216904 10338
rect 218060 4956 218112 4962
rect 218060 4898 218112 4904
rect 218072 480 218100 4898
rect 219268 480 219296 16546
rect 219452 8974 219480 79766
rect 219596 79750 219664 79778
rect 219946 79766 219998 79772
rect 220332 79778 220360 80036
rect 220694 79778 220722 80036
rect 221062 79914 221090 80036
rect 220332 79750 220400 79778
rect 219532 77308 219584 77314
rect 219532 77250 219584 77256
rect 219544 49094 219572 77250
rect 219636 49162 219664 79750
rect 220372 78130 220400 79750
rect 220648 79750 220722 79778
rect 220832 79886 221090 79914
rect 220360 78124 220412 78130
rect 220360 78066 220412 78072
rect 220648 77314 220676 79750
rect 220636 77308 220688 77314
rect 220636 77250 220688 77256
rect 219624 49156 219676 49162
rect 219624 49098 219676 49104
rect 219532 49088 219584 49094
rect 219532 49030 219584 49036
rect 219532 47592 219584 47598
rect 219532 47534 219584 47540
rect 219544 16574 219572 47534
rect 219544 16546 220032 16574
rect 219440 8968 219492 8974
rect 219440 8910 219492 8916
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220832 10538 220860 79886
rect 220912 79824 220964 79830
rect 221430 79778 221458 80036
rect 221798 79830 221826 80036
rect 220912 79766 220964 79772
rect 220924 49026 220952 79766
rect 221016 79750 221458 79778
rect 221786 79824 221838 79830
rect 221786 79766 221838 79772
rect 222172 79778 222200 80036
rect 222540 79914 222568 80036
rect 222540 79886 222608 79914
rect 222292 79824 222344 79830
rect 222172 79750 222240 79778
rect 222292 79766 222344 79772
rect 221016 56098 221044 79750
rect 221004 56092 221056 56098
rect 221004 56034 221056 56040
rect 220912 49020 220964 49026
rect 220912 48962 220964 48968
rect 222212 13258 222240 79750
rect 222304 14482 222332 79766
rect 222580 78062 222608 79886
rect 222902 79778 222930 80036
rect 223270 79830 223298 80036
rect 222856 79750 222930 79778
rect 223258 79824 223310 79830
rect 223258 79766 223310 79772
rect 223644 79778 223672 80036
rect 224006 79778 224034 80036
rect 224282 79778 224310 80036
rect 223644 79750 223712 79778
rect 222568 78056 222620 78062
rect 222568 77998 222620 78004
rect 222856 64874 222884 79750
rect 223684 77314 223712 79750
rect 223776 79750 224034 79778
rect 224236 79750 224310 79778
rect 224656 79778 224684 80036
rect 225018 79914 225046 80036
rect 224880 79886 225046 79914
rect 225386 79898 225414 80036
rect 225374 79892 225426 79898
rect 224656 79750 224724 79778
rect 223672 77308 223724 77314
rect 223672 77250 223724 77256
rect 223580 77240 223632 77246
rect 223580 77182 223632 77188
rect 222396 64846 222884 64874
rect 222396 50522 222424 64846
rect 222384 50516 222436 50522
rect 222384 50458 222436 50464
rect 222384 35284 222436 35290
rect 222384 35226 222436 35232
rect 222396 16574 222424 35226
rect 222396 16546 222792 16574
rect 222292 14476 222344 14482
rect 222292 14418 222344 14424
rect 222200 13252 222252 13258
rect 222200 13194 222252 13200
rect 220820 10532 220872 10538
rect 220820 10474 220872 10480
rect 221556 4888 221608 4894
rect 221556 4830 221608 4836
rect 221568 480 221596 4830
rect 222764 480 222792 16546
rect 223592 15910 223620 77182
rect 223672 60036 223724 60042
rect 223672 59978 223724 59984
rect 223580 15904 223632 15910
rect 223580 15846 223632 15852
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223684 354 223712 59978
rect 223776 50454 223804 79750
rect 223856 77308 223908 77314
rect 223856 77250 223908 77256
rect 223868 57458 223896 77250
rect 224236 77246 224264 79750
rect 224696 77994 224724 79750
rect 224880 79694 224908 79886
rect 225374 79834 225426 79840
rect 224960 79824 225012 79830
rect 224960 79766 225012 79772
rect 225052 79824 225104 79830
rect 225754 79778 225782 80036
rect 226122 79830 226150 80036
rect 225052 79766 225104 79772
rect 224868 79688 224920 79694
rect 224868 79630 224920 79636
rect 224684 77988 224736 77994
rect 224684 77930 224736 77936
rect 224224 77240 224276 77246
rect 224224 77182 224276 77188
rect 223856 57452 223908 57458
rect 223856 57394 223908 57400
rect 223764 50448 223816 50454
rect 223764 50390 223816 50396
rect 224972 31074 225000 79766
rect 225064 50386 225092 79766
rect 225156 79750 225782 79778
rect 226110 79824 226162 79830
rect 226490 79778 226518 80036
rect 226864 79914 226892 80036
rect 226864 79886 226932 79914
rect 226110 79766 226162 79772
rect 226352 79750 226518 79778
rect 225156 58886 225184 79750
rect 225236 79688 225288 79694
rect 225236 79630 225288 79636
rect 225248 76634 225276 79630
rect 225236 76628 225288 76634
rect 225236 76570 225288 76576
rect 225144 58880 225196 58886
rect 225144 58822 225196 58828
rect 225052 50380 225104 50386
rect 225052 50322 225104 50328
rect 224960 31068 225012 31074
rect 224960 31010 225012 31016
rect 226352 13190 226380 79750
rect 226904 78266 226932 79886
rect 227226 79778 227254 80036
rect 227594 79778 227622 80036
rect 227968 79914 227996 80036
rect 227968 79886 228036 79914
rect 227180 79750 227254 79778
rect 227548 79750 227622 79778
rect 227720 79824 227772 79830
rect 227720 79766 227772 79772
rect 226892 78260 226944 78266
rect 226892 78202 226944 78208
rect 226984 78192 227036 78198
rect 226984 78134 227036 78140
rect 226432 77308 226484 77314
rect 226432 77250 226484 77256
rect 226444 33794 226472 77250
rect 226524 77240 226576 77246
rect 226524 77182 226576 77188
rect 226536 51882 226564 77182
rect 226524 51876 226576 51882
rect 226524 51818 226576 51824
rect 226996 47870 227024 78134
rect 227180 77246 227208 79750
rect 227548 77314 227576 79750
rect 227536 77308 227588 77314
rect 227536 77250 227588 77256
rect 227168 77240 227220 77246
rect 227168 77182 227220 77188
rect 226984 47864 227036 47870
rect 226984 47806 227036 47812
rect 226524 42084 226576 42090
rect 226524 42026 226576 42032
rect 226432 33788 226484 33794
rect 226432 33730 226484 33736
rect 226340 13184 226392 13190
rect 226340 13126 226392 13132
rect 226536 6914 226564 42026
rect 227732 10470 227760 79766
rect 228008 78334 228036 79886
rect 228330 79778 228358 80036
rect 228698 79830 228726 80036
rect 229066 79914 229094 80036
rect 229066 79886 229232 79914
rect 228100 79750 228358 79778
rect 228686 79824 228738 79830
rect 228686 79766 228738 79772
rect 229100 79824 229152 79830
rect 229100 79766 229152 79772
rect 227996 78328 228048 78334
rect 227996 78270 228048 78276
rect 228100 64874 228128 79750
rect 227824 64846 228128 64874
rect 227824 22846 227852 64846
rect 227812 22840 227864 22846
rect 227812 22782 227864 22788
rect 227720 10464 227772 10470
rect 227720 10406 227772 10412
rect 229112 10402 229140 79766
rect 229204 77450 229232 79886
rect 229434 79778 229462 80036
rect 229802 79898 229830 80036
rect 229790 79892 229842 79898
rect 229790 79834 229842 79840
rect 230170 79778 230198 80036
rect 229388 79750 229462 79778
rect 229664 79750 230198 79778
rect 230544 79778 230572 80036
rect 230906 79898 230934 80036
rect 231274 79898 231302 80036
rect 230894 79892 230946 79898
rect 230894 79834 230946 79840
rect 231262 79892 231314 79898
rect 231262 79834 231314 79840
rect 231642 79778 231670 80036
rect 231860 79892 231912 79898
rect 231860 79834 231912 79840
rect 230544 79750 230704 79778
rect 229192 77444 229244 77450
rect 229192 77386 229244 77392
rect 229388 77330 229416 79750
rect 229204 77302 229416 77330
rect 229204 42090 229232 77302
rect 229284 77240 229336 77246
rect 229284 77182 229336 77188
rect 229296 44878 229324 77182
rect 229664 64874 229692 79750
rect 230480 79688 230532 79694
rect 230480 79630 230532 79636
rect 230572 79688 230624 79694
rect 230572 79630 230624 79636
rect 229388 64846 229692 64874
rect 229388 61402 229416 64846
rect 229376 61396 229428 61402
rect 229376 61338 229428 61344
rect 229284 44872 229336 44878
rect 229284 44814 229336 44820
rect 229192 42084 229244 42090
rect 229192 42026 229244 42032
rect 229192 26920 229244 26926
rect 229192 26862 229244 26868
rect 229204 16574 229232 26862
rect 229204 16546 229416 16574
rect 229100 10396 229152 10402
rect 229100 10338 229152 10344
rect 227536 10328 227588 10334
rect 227536 10270 227588 10276
rect 226352 6886 226564 6914
rect 225144 5160 225196 5166
rect 225144 5102 225196 5108
rect 225156 480 225184 5102
rect 226352 480 226380 6886
rect 227548 480 227576 10270
rect 228732 4820 228784 4826
rect 228732 4762 228784 4768
rect 228744 480 228772 4762
rect 223918 354 224030 480
rect 223684 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 16546
rect 230492 10334 230520 79630
rect 230584 11966 230612 79630
rect 230676 24342 230704 79750
rect 230768 79750 231670 79778
rect 230664 24336 230716 24342
rect 230664 24278 230716 24284
rect 230768 24274 230796 79750
rect 230756 24268 230808 24274
rect 230756 24210 230808 24216
rect 231872 17474 231900 79834
rect 232016 79778 232044 80036
rect 232378 79898 232406 80036
rect 232746 79898 232774 80036
rect 232366 79892 232418 79898
rect 232366 79834 232418 79840
rect 232734 79892 232786 79898
rect 232734 79834 232786 79840
rect 233114 79778 233142 80036
rect 233482 79778 233510 80036
rect 233850 79778 233878 80036
rect 234218 79778 234246 80036
rect 232016 79750 232084 79778
rect 231952 79688 232004 79694
rect 231952 79630 232004 79636
rect 231964 24206 231992 79630
rect 232056 51814 232084 79750
rect 232148 79750 233142 79778
rect 233252 79750 233510 79778
rect 233620 79750 233878 79778
rect 234172 79750 234246 79778
rect 234592 79778 234620 80036
rect 234954 79778 234982 80036
rect 235322 79778 235350 80036
rect 235690 79778 235718 80036
rect 234592 79750 234752 79778
rect 232044 51808 232096 51814
rect 232044 51750 232096 51756
rect 232148 51746 232176 79750
rect 232136 51740 232188 51746
rect 232136 51682 232188 51688
rect 231952 24200 232004 24206
rect 231952 24142 232004 24148
rect 231952 18692 232004 18698
rect 231952 18634 232004 18640
rect 231860 17468 231912 17474
rect 231860 17410 231912 17416
rect 230572 11960 230624 11966
rect 230572 11902 230624 11908
rect 231032 10668 231084 10674
rect 231032 10610 231084 10616
rect 230480 10328 230532 10334
rect 230480 10270 230532 10276
rect 231044 480 231072 10610
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231964 354 231992 18634
rect 233252 17406 233280 79750
rect 233620 77330 233648 79750
rect 233344 77302 233648 77330
rect 233344 25702 233372 77302
rect 234172 64874 234200 79750
rect 234620 77308 234672 77314
rect 234620 77250 234672 77256
rect 233436 64846 234200 64874
rect 233436 53242 233464 64846
rect 233424 53236 233476 53242
rect 233424 53178 233476 53184
rect 233424 35216 233476 35222
rect 233424 35158 233476 35164
rect 233332 25696 233384 25702
rect 233332 25638 233384 25644
rect 233240 17400 233292 17406
rect 233240 17342 233292 17348
rect 233436 480 233464 35158
rect 234632 17270 234660 77250
rect 234724 17338 234752 79750
rect 234816 79750 234982 79778
rect 235276 79750 235350 79778
rect 235644 79750 235718 79778
rect 236064 79778 236092 80036
rect 236334 79778 236362 80036
rect 236702 79778 236730 80036
rect 237070 79778 237098 80036
rect 236064 79750 236224 79778
rect 234816 25634 234844 79750
rect 235276 64874 235304 79750
rect 235644 77314 235672 79750
rect 235632 77308 235684 77314
rect 235632 77250 235684 77256
rect 236092 77308 236144 77314
rect 236092 77250 236144 77256
rect 236000 77240 236052 77246
rect 236000 77182 236052 77188
rect 234908 64846 235304 64874
rect 234908 53174 234936 64846
rect 234896 53168 234948 53174
rect 234896 53110 234948 53116
rect 234896 50720 234948 50726
rect 234896 50662 234948 50668
rect 234804 25628 234856 25634
rect 234804 25570 234856 25576
rect 234804 18624 234856 18630
rect 234804 18566 234856 18572
rect 234712 17332 234764 17338
rect 234712 17274 234764 17280
rect 234620 17264 234672 17270
rect 234620 17206 234672 17212
rect 234816 12782 234844 18566
rect 234804 12776 234856 12782
rect 234804 12718 234856 12724
rect 234908 6914 234936 50662
rect 236012 25566 236040 77182
rect 236104 36582 236132 77250
rect 236196 43450 236224 79750
rect 236288 79750 236362 79778
rect 236656 79750 236730 79778
rect 237024 79750 237098 79778
rect 237444 79778 237472 80036
rect 237806 79778 237834 80036
rect 238174 79898 238202 80036
rect 238162 79892 238214 79898
rect 238162 79834 238214 79840
rect 238542 79778 238570 80036
rect 237444 79750 237512 79778
rect 236288 53106 236316 79750
rect 236656 77314 236684 79750
rect 236644 77308 236696 77314
rect 236644 77250 236696 77256
rect 237024 77246 237052 79750
rect 237380 79688 237432 79694
rect 237380 79630 237432 79636
rect 237012 77240 237064 77246
rect 237012 77182 237064 77188
rect 236276 53100 236328 53106
rect 236276 53042 236328 53048
rect 236184 43444 236236 43450
rect 236184 43386 236236 43392
rect 236184 36916 236236 36922
rect 236184 36858 236236 36864
rect 236092 36576 236144 36582
rect 236092 36518 236144 36524
rect 236000 25560 236052 25566
rect 236000 25502 236052 25508
rect 236196 16574 236224 36858
rect 237392 27062 237420 79630
rect 237484 54738 237512 79750
rect 237576 79750 237834 79778
rect 237944 79750 238570 79778
rect 238760 79824 238812 79830
rect 238910 79778 238938 80036
rect 239278 79778 239306 80036
rect 239646 79830 239674 80036
rect 238760 79766 238812 79772
rect 237472 54732 237524 54738
rect 237472 54674 237524 54680
rect 237472 52080 237524 52086
rect 237472 52022 237524 52028
rect 237380 27056 237432 27062
rect 237380 26998 237432 27004
rect 237484 16574 237512 52022
rect 237576 37942 237604 79750
rect 237944 64874 237972 79750
rect 237668 64846 237972 64874
rect 237668 54670 237696 64846
rect 237656 54664 237708 54670
rect 237656 54606 237708 54612
rect 238772 54602 238800 79766
rect 238864 79750 238938 79778
rect 239048 79750 239306 79778
rect 239634 79824 239686 79830
rect 240014 79778 240042 80036
rect 240382 79880 240410 80036
rect 239634 79766 239686 79772
rect 239968 79750 240042 79778
rect 240152 79852 240410 79880
rect 238864 62830 238892 79750
rect 238944 77308 238996 77314
rect 238944 77250 238996 77256
rect 238956 64190 238984 77250
rect 239048 73982 239076 79750
rect 239968 77314 239996 79750
rect 239956 77308 240008 77314
rect 239956 77250 240008 77256
rect 239036 73976 239088 73982
rect 239036 73918 239088 73924
rect 238944 64184 238996 64190
rect 238944 64126 238996 64132
rect 238852 62824 238904 62830
rect 238852 62766 238904 62772
rect 238760 54596 238812 54602
rect 238760 54538 238812 54544
rect 237564 37936 237616 37942
rect 237564 37878 237616 37884
rect 238760 18828 238812 18834
rect 238760 18770 238812 18776
rect 238772 16574 238800 18770
rect 236196 16546 236592 16574
rect 237484 16546 237696 16574
rect 238772 16546 239352 16574
rect 235816 12776 235868 12782
rect 235816 12718 235868 12724
rect 234632 6886 234936 6914
rect 234632 480 234660 6886
rect 235828 480 235856 12718
rect 232198 354 232310 480
rect 231964 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 240152 4962 240180 79852
rect 240750 79778 240778 80036
rect 241118 79778 241146 80036
rect 240336 79750 240778 79778
rect 241072 79750 241146 79778
rect 241492 79778 241520 80036
rect 241704 79824 241756 79830
rect 241492 79750 241652 79778
rect 241854 79778 241882 80036
rect 242222 79778 242250 80036
rect 242590 79830 242618 80036
rect 241704 79766 241756 79772
rect 240232 77308 240284 77314
rect 240232 77250 240284 77256
rect 240244 22778 240272 77250
rect 240336 56030 240364 79750
rect 241072 77314 241100 79750
rect 241060 77308 241112 77314
rect 241060 77250 241112 77256
rect 241520 77308 241572 77314
rect 241520 77250 241572 77256
rect 240324 56024 240376 56030
rect 240324 55966 240376 55972
rect 240324 38276 240376 38282
rect 240324 38218 240376 38224
rect 240232 22772 240284 22778
rect 240232 22714 240284 22720
rect 240140 4956 240192 4962
rect 240140 4898 240192 4904
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240336 354 240364 38218
rect 241532 24138 241560 77250
rect 241624 26994 241652 79750
rect 241612 26988 241664 26994
rect 241612 26930 241664 26936
rect 241716 26926 241744 79766
rect 241808 79750 241882 79778
rect 242176 79750 242250 79778
rect 242578 79824 242630 79830
rect 242578 79766 242630 79772
rect 242964 79778 242992 80036
rect 243326 79778 243354 80036
rect 243694 79778 243722 80036
rect 244062 79778 244090 80036
rect 244280 79892 244332 79898
rect 244280 79834 244332 79840
rect 242964 79750 243216 79778
rect 241808 55962 241836 79750
rect 242176 77314 242204 79750
rect 242992 77376 243044 77382
rect 242992 77318 243044 77324
rect 242164 77308 242216 77314
rect 242164 77250 242216 77256
rect 242900 77240 242952 77246
rect 242900 77182 242952 77188
rect 241796 55956 241848 55962
rect 241796 55898 241848 55904
rect 242912 40798 242940 77182
rect 243004 55894 243032 77318
rect 243084 77308 243136 77314
rect 243084 77250 243136 77256
rect 243096 72554 243124 77250
rect 243188 73914 243216 79750
rect 243280 79750 243354 79778
rect 243648 79750 243722 79778
rect 244016 79750 244090 79778
rect 243280 77246 243308 79750
rect 243648 77314 243676 79750
rect 244016 77382 244044 79750
rect 244004 77376 244056 77382
rect 244004 77318 244056 77324
rect 243636 77308 243688 77314
rect 243636 77250 243688 77256
rect 243268 77240 243320 77246
rect 243268 77182 243320 77188
rect 243176 73908 243228 73914
rect 243176 73850 243228 73856
rect 243084 72548 243136 72554
rect 243084 72490 243136 72496
rect 242992 55888 243044 55894
rect 242992 55830 243044 55836
rect 242900 40792 242952 40798
rect 242900 40734 242952 40740
rect 242900 39364 242952 39370
rect 242900 39306 242952 39312
rect 241704 26920 241756 26926
rect 241704 26862 241756 26868
rect 241520 24132 241572 24138
rect 241520 24074 241572 24080
rect 241704 11892 241756 11898
rect 241704 11834 241756 11840
rect 241716 480 241744 11834
rect 242912 11830 242940 39306
rect 244292 28422 244320 79834
rect 244430 79778 244458 80036
rect 244798 79898 244826 80036
rect 244786 79892 244838 79898
rect 244786 79834 244838 79840
rect 245166 79778 245194 80036
rect 245534 79778 245562 80036
rect 245902 79880 245930 80036
rect 244384 79750 244458 79778
rect 244568 79750 245194 79778
rect 245488 79750 245562 79778
rect 245672 79852 245930 79880
rect 244384 39370 244412 79750
rect 244464 77308 244516 77314
rect 244464 77250 244516 77256
rect 244476 47598 244504 77250
rect 244568 57390 244596 79750
rect 245488 77314 245516 79750
rect 245476 77308 245528 77314
rect 245476 77250 245528 77256
rect 244556 57384 244608 57390
rect 244556 57326 244608 57332
rect 244464 47592 244516 47598
rect 244464 47534 244516 47540
rect 244372 39364 244424 39370
rect 244372 39306 244424 39312
rect 244280 28416 244332 28422
rect 244280 28358 244332 28364
rect 242992 24540 243044 24546
rect 242992 24482 243044 24488
rect 242900 11824 242952 11830
rect 242900 11766 242952 11772
rect 243004 6914 243032 24482
rect 245200 11892 245252 11898
rect 245200 11834 245252 11840
rect 244096 11824 244148 11830
rect 244096 11766 244148 11772
rect 242912 6886 243032 6914
rect 242912 480 242940 6886
rect 244108 480 244136 11766
rect 245212 480 245240 11834
rect 245672 4894 245700 79852
rect 246270 79778 246298 80036
rect 246638 79778 246666 80036
rect 245856 79750 246298 79778
rect 246592 79750 246666 79778
rect 247012 79778 247040 80036
rect 247374 79778 247402 80036
rect 247742 79778 247770 80036
rect 248110 79778 248138 80036
rect 248392 79914 248420 80036
rect 248392 79886 248644 79914
rect 248760 79898 248788 80036
rect 247012 79750 247264 79778
rect 245752 77308 245804 77314
rect 245752 77250 245804 77256
rect 245764 18834 245792 77250
rect 245856 57322 245884 79750
rect 246592 77314 246620 79750
rect 246580 77308 246632 77314
rect 246580 77250 246632 77256
rect 247132 77308 247184 77314
rect 247132 77250 247184 77256
rect 247040 77240 247092 77246
rect 247040 77182 247092 77188
rect 247052 60110 247080 77182
rect 247144 65550 247172 77250
rect 247236 72486 247264 79750
rect 247328 79750 247402 79778
rect 247696 79750 247770 79778
rect 248064 79750 248138 79778
rect 248420 79824 248472 79830
rect 248420 79766 248472 79772
rect 247328 73846 247356 79750
rect 247696 77314 247724 79750
rect 247684 77308 247736 77314
rect 247684 77250 247736 77256
rect 248064 77246 248092 79750
rect 248052 77240 248104 77246
rect 248052 77182 248104 77188
rect 247316 73840 247368 73846
rect 247316 73782 247368 73788
rect 247224 72480 247276 72486
rect 247224 72422 247276 72428
rect 247132 65544 247184 65550
rect 247132 65486 247184 65492
rect 247040 60104 247092 60110
rect 247040 60046 247092 60052
rect 245844 57316 245896 57322
rect 245844 57258 245896 57264
rect 247040 43784 247092 43790
rect 247040 43726 247092 43732
rect 245844 24472 245896 24478
rect 245844 24414 245896 24420
rect 245752 18828 245804 18834
rect 245752 18770 245804 18776
rect 245856 16574 245884 24414
rect 247052 16574 247080 43726
rect 245856 16546 245976 16574
rect 247052 16546 247632 16574
rect 245660 4888 245712 4894
rect 245660 4830 245712 4836
rect 240478 354 240590 480
rect 240336 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 248432 4826 248460 79766
rect 248512 77308 248564 77314
rect 248512 77250 248564 77256
rect 248524 11898 248552 77250
rect 248616 57254 248644 79886
rect 248748 79892 248800 79898
rect 248748 79834 248800 79840
rect 249122 79830 249150 80036
rect 249110 79824 249162 79830
rect 249490 79778 249518 80036
rect 249616 79892 249668 79898
rect 249616 79834 249668 79840
rect 249110 79766 249162 79772
rect 249444 79750 249518 79778
rect 249444 77314 249472 79750
rect 249432 77308 249484 77314
rect 249432 77250 249484 77256
rect 249628 75206 249656 79834
rect 249864 79778 249892 80036
rect 250226 79778 250254 80036
rect 250594 79914 250622 80036
rect 249864 79750 249932 79778
rect 249800 77308 249852 77314
rect 249800 77250 249852 77256
rect 249616 75200 249668 75206
rect 249616 75142 249668 75148
rect 248604 57248 248656 57254
rect 248604 57190 248656 57196
rect 248512 11892 248564 11898
rect 248512 11834 248564 11840
rect 249812 11830 249840 77250
rect 249904 13122 249932 79750
rect 249996 79750 250254 79778
rect 250364 79886 250622 79914
rect 249996 28354 250024 79750
rect 250364 77314 250392 79886
rect 250962 79778 250990 80036
rect 251180 79892 251232 79898
rect 251180 79834 251232 79840
rect 250456 79750 250990 79778
rect 250352 77308 250404 77314
rect 250352 77250 250404 77256
rect 250456 66910 250484 79750
rect 250444 66904 250496 66910
rect 250444 66846 250496 66852
rect 249984 28348 250036 28354
rect 249984 28290 250036 28296
rect 249984 25900 250036 25906
rect 249984 25842 250036 25848
rect 249892 13116 249944 13122
rect 249892 13058 249944 13064
rect 249800 11824 249852 11830
rect 249800 11766 249852 11772
rect 248512 11756 248564 11762
rect 248512 11698 248564 11704
rect 248420 4820 248472 4826
rect 248420 4762 248472 4768
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248524 354 248552 11698
rect 249996 480 250024 25842
rect 251192 11762 251220 79834
rect 251330 79778 251358 80036
rect 251698 79898 251726 80036
rect 251686 79892 251738 79898
rect 251686 79834 251738 79840
rect 252066 79778 252094 80036
rect 252434 79778 252462 80036
rect 252652 79892 252704 79898
rect 252652 79834 252704 79840
rect 251284 79750 251358 79778
rect 251468 79750 252094 79778
rect 252388 79750 252462 79778
rect 252560 79824 252612 79830
rect 252560 79766 252612 79772
rect 251284 28286 251312 79750
rect 251364 77308 251416 77314
rect 251364 77250 251416 77256
rect 251376 29782 251404 77250
rect 251468 68338 251496 79750
rect 252388 77314 252416 79750
rect 252376 77308 252428 77314
rect 252376 77250 252428 77256
rect 251456 68332 251508 68338
rect 251456 68274 251508 68280
rect 251456 46504 251508 46510
rect 251456 46446 251508 46452
rect 251364 29776 251416 29782
rect 251364 29718 251416 29724
rect 251272 28280 251324 28286
rect 251272 28222 251324 28228
rect 251272 13456 251324 13462
rect 251272 13398 251324 13404
rect 251180 11756 251232 11762
rect 251180 11698 251232 11704
rect 251284 3602 251312 13398
rect 251468 6914 251496 46446
rect 252572 18766 252600 79766
rect 252664 29714 252692 79834
rect 252802 79778 252830 80036
rect 253170 79830 253198 80036
rect 253538 79898 253566 80036
rect 253526 79892 253578 79898
rect 253526 79834 253578 79840
rect 252756 79750 252830 79778
rect 253158 79824 253210 79830
rect 253158 79766 253210 79772
rect 253912 79778 253940 80036
rect 254124 79892 254176 79898
rect 254124 79834 254176 79840
rect 254032 79824 254084 79830
rect 253912 79750 253980 79778
rect 254032 79766 254084 79772
rect 252756 40730 252784 79750
rect 253952 58818 253980 79750
rect 253940 58812 253992 58818
rect 253940 58754 253992 58760
rect 253940 47932 253992 47938
rect 253940 47874 253992 47880
rect 252744 40724 252796 40730
rect 252744 40666 252796 40672
rect 252652 29708 252704 29714
rect 252652 29650 252704 29656
rect 252652 25832 252704 25838
rect 252652 25774 252704 25780
rect 252560 18760 252612 18766
rect 252560 18702 252612 18708
rect 252664 16574 252692 25774
rect 253952 16574 253980 47874
rect 254044 35358 254072 79766
rect 254136 58750 254164 79834
rect 254274 79778 254302 80036
rect 254642 79830 254670 80036
rect 255010 79898 255038 80036
rect 254998 79892 255050 79898
rect 254998 79834 255050 79840
rect 254228 79750 254302 79778
rect 254630 79824 254682 79830
rect 255378 79778 255406 80036
rect 255746 79778 255774 80036
rect 256114 79778 256142 80036
rect 256482 79778 256510 80036
rect 256850 79914 256878 80036
rect 254630 79766 254682 79772
rect 255332 79750 255406 79778
rect 255516 79750 255774 79778
rect 255884 79750 256142 79778
rect 256436 79750 256510 79778
rect 256712 79886 256878 79914
rect 254228 69698 254256 79750
rect 254216 69692 254268 69698
rect 254216 69634 254268 69640
rect 254124 58744 254176 58750
rect 254124 58686 254176 58692
rect 254032 35352 254084 35358
rect 254032 35294 254084 35300
rect 255332 18698 255360 79750
rect 255516 77330 255544 79750
rect 255424 77302 255544 77330
rect 255424 29646 255452 77302
rect 255884 77194 255912 79750
rect 255964 78124 256016 78130
rect 255964 78066 256016 78072
rect 255516 77166 255912 77194
rect 255516 58682 255544 77166
rect 255596 77104 255648 77110
rect 255596 77046 255648 77052
rect 255608 71058 255636 77046
rect 255596 71052 255648 71058
rect 255596 70994 255648 71000
rect 255504 58676 255556 58682
rect 255504 58618 255556 58624
rect 255412 29640 255464 29646
rect 255412 29582 255464 29588
rect 255320 18692 255372 18698
rect 255320 18634 255372 18640
rect 252664 16546 253520 16574
rect 253952 16546 254256 16574
rect 251376 6886 251496 6914
rect 251272 3596 251324 3602
rect 251272 3538 251324 3544
rect 251376 3482 251404 6886
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 251192 3454 251404 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3538
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248524 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255976 13326 256004 78066
rect 256436 77110 256464 79750
rect 256424 77104 256476 77110
rect 256424 77046 256476 77052
rect 256712 35290 256740 79886
rect 256792 79824 256844 79830
rect 257218 79778 257246 80036
rect 256792 79766 256844 79772
rect 256700 35284 256752 35290
rect 256700 35226 256752 35232
rect 256804 35222 256832 79766
rect 256896 79750 257246 79778
rect 257592 79778 257620 80036
rect 257954 79830 257982 80036
rect 257942 79824 257994 79830
rect 257592 79750 257660 79778
rect 257942 79766 257994 79772
rect 258080 79824 258132 79830
rect 258322 79778 258350 80036
rect 258690 79830 258718 80036
rect 258080 79766 258132 79772
rect 256896 54534 256924 79750
rect 257632 76566 257660 79750
rect 257620 76560 257672 76566
rect 257620 76502 257672 76508
rect 256884 54528 256936 54534
rect 256884 54470 256936 54476
rect 256792 35216 256844 35222
rect 256792 35158 256844 35164
rect 256700 22976 256752 22982
rect 256700 22918 256752 22924
rect 255872 13320 255924 13326
rect 255872 13262 255924 13268
rect 255964 13320 256016 13326
rect 255964 13262 256016 13268
rect 255884 480 255912 13262
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 22918
rect 258092 18630 258120 79766
rect 258184 79750 258350 79778
rect 258678 79824 258730 79830
rect 258678 79766 258730 79772
rect 259064 79778 259092 80036
rect 259432 79778 259460 80036
rect 259808 80022 260144 80050
rect 259064 79750 259132 79778
rect 259432 79750 259500 79778
rect 258184 60042 258212 79750
rect 258724 78328 258776 78334
rect 258724 78270 258776 78276
rect 258172 60036 258224 60042
rect 258172 59978 258224 59984
rect 258172 49292 258224 49298
rect 258172 49234 258224 49240
rect 258080 18624 258132 18630
rect 258080 18566 258132 18572
rect 258184 16574 258212 49234
rect 258184 16546 258304 16574
rect 258276 480 258304 16546
rect 258736 3670 258764 78270
rect 259104 78198 259132 79750
rect 259092 78192 259144 78198
rect 259092 78134 259144 78140
rect 258724 3664 258776 3670
rect 258724 3606 258776 3612
rect 259472 3602 259500 79750
rect 260116 78130 260144 80022
rect 260104 78124 260156 78130
rect 260104 78066 260156 78072
rect 259552 64456 259604 64462
rect 259552 64398 259604 64404
rect 259460 3596 259512 3602
rect 259460 3538 259512 3544
rect 259564 3482 259592 64398
rect 260840 50652 260892 50658
rect 260840 50594 260892 50600
rect 259644 27260 259696 27266
rect 259644 27202 259696 27208
rect 259656 16574 259684 27202
rect 260852 16574 260880 50594
rect 261496 46918 261524 200466
rect 261588 167006 261616 201622
rect 445496 200802 445524 419834
rect 445588 200938 445616 419999
rect 520660 419914 520688 421126
rect 520414 419886 520688 419914
rect 445668 419824 445720 419830
rect 521028 419778 521056 421262
rect 521568 421252 521620 421258
rect 521568 421194 521620 421200
rect 521198 420472 521254 420481
rect 521198 420407 521254 420416
rect 521212 419914 521240 420407
rect 521580 419914 521608 421194
rect 522040 419914 522068 422758
rect 522764 421116 522816 421122
rect 522764 421058 522816 421064
rect 522394 420472 522450 420481
rect 522394 420407 522450 420416
rect 522408 419914 522436 420407
rect 522776 419914 522804 421058
rect 522960 419914 522988 422826
rect 523776 422340 523828 422346
rect 523776 422282 523828 422288
rect 523498 421016 523554 421025
rect 523498 420951 523554 420960
rect 523512 419914 523540 420951
rect 523788 419914 523816 422282
rect 524156 419914 524184 423098
rect 529020 422748 529072 422754
rect 529020 422690 529072 422696
rect 525708 422476 525760 422482
rect 525708 422418 525760 422424
rect 525614 421152 525670 421161
rect 525614 421087 525670 421096
rect 524880 421048 524932 421054
rect 524880 420990 524932 420996
rect 524512 420436 524564 420442
rect 524512 420378 524564 420384
rect 524524 419914 524552 420378
rect 524892 419914 524920 420990
rect 525248 420980 525300 420986
rect 525248 420922 525300 420928
rect 525260 419914 525288 420922
rect 525628 419914 525656 421087
rect 525720 420186 525748 422418
rect 526260 422408 526312 422414
rect 526260 422350 526312 422356
rect 527086 422376 527142 422385
rect 525892 420504 525944 420510
rect 525892 420446 525944 420452
rect 525720 420158 525840 420186
rect 525812 419914 525840 420158
rect 521150 419886 521240 419914
rect 521518 419886 521608 419914
rect 521886 419886 522068 419914
rect 522162 419886 522436 419914
rect 522530 419886 522804 419914
rect 522898 419886 522988 419914
rect 523266 419886 523540 419914
rect 523634 419886 523816 419914
rect 523910 419886 524184 419914
rect 524278 419886 524552 419914
rect 524646 419886 524920 419914
rect 525014 419886 525288 419914
rect 525382 419886 525656 419914
rect 525750 419886 525840 419914
rect 525904 419830 525932 420446
rect 526272 419914 526300 422350
rect 527086 422311 527142 422320
rect 527100 421666 527128 422311
rect 527640 421864 527692 421870
rect 527640 421806 527692 421812
rect 527088 421660 527140 421666
rect 527088 421602 527140 421608
rect 526904 421388 526956 421394
rect 526904 421330 526956 421336
rect 526626 421288 526682 421297
rect 526626 421223 526682 421232
rect 526640 419914 526668 421223
rect 526916 419914 526944 421330
rect 527364 420028 527416 420034
rect 527364 419970 527416 419976
rect 527376 419914 527404 419970
rect 527652 419914 527680 421806
rect 528468 421796 528520 421802
rect 528468 421738 528520 421744
rect 528008 421456 528060 421462
rect 528008 421398 528060 421404
rect 528020 419914 528048 421398
rect 528480 420186 528508 421738
rect 528928 421524 528980 421530
rect 528928 421466 528980 421472
rect 528480 420158 528600 420186
rect 528572 419914 528600 420158
rect 528940 419914 528968 421466
rect 526026 419886 526300 419914
rect 526394 419886 526668 419914
rect 526762 419886 526944 419914
rect 527130 419886 527404 419914
rect 527498 419886 527680 419914
rect 527774 419886 528048 419914
rect 528510 419886 528600 419914
rect 528878 419886 528968 419914
rect 445668 419766 445720 419772
rect 445576 200932 445628 200938
rect 445576 200874 445628 200880
rect 445680 200870 445708 419766
rect 520782 419750 521056 419778
rect 525892 419824 525944 419830
rect 528376 419824 528428 419830
rect 525892 419766 525944 419772
rect 528142 419772 528376 419778
rect 528142 419766 528428 419772
rect 529032 419778 529060 422690
rect 529216 420918 529244 424322
rect 529296 421932 529348 421938
rect 529296 421874 529348 421880
rect 529204 420912 529256 420918
rect 529204 420854 529256 420860
rect 529308 419914 529336 421874
rect 529480 420096 529532 420102
rect 529480 420038 529532 420044
rect 529492 419914 529520 420038
rect 529676 419914 529704 430578
rect 530136 423638 530164 484366
rect 530584 456816 530636 456822
rect 530584 456758 530636 456764
rect 530596 441614 530624 456758
rect 530596 441586 530808 441614
rect 530124 423632 530176 423638
rect 530124 423574 530176 423580
rect 530492 422612 530544 422618
rect 530492 422554 530544 422560
rect 529940 422340 529992 422346
rect 529940 422282 529992 422288
rect 529952 421666 529980 422282
rect 529940 421660 529992 421666
rect 529940 421602 529992 421608
rect 530124 420368 530176 420374
rect 530124 420310 530176 420316
rect 530032 420300 530084 420306
rect 530032 420242 530084 420248
rect 530044 419966 530072 420242
rect 530032 419960 530084 419966
rect 529308 419886 529598 419914
rect 529676 419886 529874 419914
rect 530032 419902 530084 419908
rect 530136 419898 530164 420310
rect 530504 419914 530532 422554
rect 530780 422006 530808 441586
rect 531332 423638 531360 524418
rect 531412 470620 531464 470626
rect 531412 470562 531464 470568
rect 530860 423632 530912 423638
rect 530860 423574 530912 423580
rect 531320 423632 531372 423638
rect 531320 423574 531372 423580
rect 530768 422000 530820 422006
rect 530768 421942 530820 421948
rect 530124 419892 530176 419898
rect 530258 419886 530532 419914
rect 530124 419834 530176 419840
rect 530780 419778 530808 421942
rect 530872 419914 530900 423574
rect 531424 419914 531452 470562
rect 531872 427440 531924 427446
rect 531872 427382 531924 427388
rect 531688 424448 531740 424454
rect 531688 424390 531740 424396
rect 531700 420170 531728 424390
rect 531688 420164 531740 420170
rect 531688 420106 531740 420112
rect 531700 419914 531728 420106
rect 530872 419886 530978 419914
rect 531362 419886 531452 419914
rect 531638 419886 531728 419914
rect 531884 419914 531912 427382
rect 532804 424726 532832 576846
rect 532792 424720 532844 424726
rect 532792 424662 532844 424668
rect 532792 424516 532844 424522
rect 532792 424458 532844 424464
rect 532056 423632 532108 423638
rect 532056 423574 532108 423580
rect 532068 419914 532096 423574
rect 532804 421734 532832 424458
rect 532792 421728 532844 421734
rect 532792 421670 532844 421676
rect 532804 419914 532832 421670
rect 531884 419886 531990 419914
rect 532068 419886 532358 419914
rect 532742 419886 532832 419914
rect 532896 419914 532924 590650
rect 533356 427814 533384 616830
rect 534184 427814 534212 630634
rect 534368 441614 534396 696934
rect 535552 683188 535604 683194
rect 535552 683130 535604 683136
rect 534368 441586 534948 441614
rect 533356 427786 533568 427814
rect 534184 427786 534580 427814
rect 533160 424720 533212 424726
rect 533160 424662 533212 424668
rect 533172 419914 533200 424662
rect 533540 423298 533568 427786
rect 534356 427508 534408 427514
rect 534356 427450 534408 427456
rect 533528 423292 533580 423298
rect 533528 423234 533580 423240
rect 533540 419914 533568 423234
rect 532896 419886 533094 419914
rect 533172 419886 533462 419914
rect 533540 419886 533738 419914
rect 534368 419778 534396 427450
rect 534552 419914 534580 427786
rect 534724 422680 534776 422686
rect 534724 422622 534776 422628
rect 534490 419886 534580 419914
rect 534736 419914 534764 422622
rect 534920 419914 534948 441586
rect 535184 425944 535236 425950
rect 535184 425886 535236 425892
rect 535196 422686 535224 425886
rect 535184 422680 535236 422686
rect 535184 422622 535236 422628
rect 535276 422680 535328 422686
rect 535276 422622 535328 422628
rect 535288 421841 535316 422622
rect 535368 422476 535420 422482
rect 535368 422418 535420 422424
rect 535274 421832 535330 421841
rect 535274 421767 535330 421776
rect 535380 421734 535408 422418
rect 535368 421728 535420 421734
rect 535368 421670 535420 421676
rect 535564 419914 535592 683130
rect 535644 453348 535696 453354
rect 535644 453290 535696 453296
rect 535656 427814 535684 453290
rect 535748 441614 535776 700470
rect 543004 700460 543056 700466
rect 543004 700402 543056 700408
rect 542636 599616 542688 599622
rect 542636 599558 542688 599564
rect 539876 510672 539928 510678
rect 539876 510614 539928 510620
rect 536840 497548 536892 497554
rect 536840 497490 536892 497496
rect 536852 441614 536880 497490
rect 539692 497480 539744 497486
rect 539692 497422 539744 497428
rect 535748 441586 536328 441614
rect 536852 441586 537340 441614
rect 535656 427786 535960 427814
rect 535736 423224 535788 423230
rect 535736 423166 535788 423172
rect 534736 419886 534842 419914
rect 534920 419886 535210 419914
rect 535502 419886 535592 419914
rect 535748 419914 535776 423166
rect 535932 419914 535960 427786
rect 536300 419914 536328 441586
rect 537024 427372 537076 427378
rect 537024 427314 537076 427320
rect 536840 424652 536892 424658
rect 536840 424594 536892 424600
rect 536748 424584 536800 424590
rect 536748 424526 536800 424532
rect 536760 423230 536788 424526
rect 536748 423224 536800 423230
rect 536748 423166 536800 423172
rect 536852 419914 536880 424594
rect 537036 419914 537064 427314
rect 537312 419914 537340 441586
rect 538496 428800 538548 428806
rect 538496 428742 538548 428748
rect 538220 427304 538272 427310
rect 538220 427246 538272 427252
rect 537668 420912 537720 420918
rect 537668 420854 537720 420860
rect 537680 419914 537708 420854
rect 538232 419914 538260 427246
rect 538508 419914 538536 428742
rect 539704 428670 539732 497422
rect 539784 428868 539836 428874
rect 539784 428810 539836 428816
rect 539692 428664 539744 428670
rect 539692 428606 539744 428612
rect 539140 425876 539192 425882
rect 539140 425818 539192 425824
rect 538864 425264 538916 425270
rect 538864 425206 538916 425212
rect 538772 422408 538824 422414
rect 538772 422350 538824 422356
rect 538784 420646 538812 422350
rect 538772 420640 538824 420646
rect 538772 420582 538824 420588
rect 538876 419914 538904 425206
rect 539152 419914 539180 425818
rect 539416 420504 539468 420510
rect 539416 420446 539468 420452
rect 539428 420170 539456 420446
rect 539416 420164 539468 420170
rect 539416 420106 539468 420112
rect 539796 419914 539824 428810
rect 535748 419886 535854 419914
rect 535932 419886 536222 419914
rect 536300 419886 536590 419914
rect 536852 419886 536958 419914
rect 537036 419886 537234 419914
rect 537312 419886 537602 419914
rect 537680 419886 537970 419914
rect 538232 419886 538338 419914
rect 538508 419886 538706 419914
rect 538876 419886 539074 419914
rect 539152 419886 539350 419914
rect 539734 419886 539824 419914
rect 539888 419914 539916 510614
rect 541532 428800 541584 428806
rect 541532 428742 541584 428748
rect 540520 428664 540572 428670
rect 540520 428606 540572 428612
rect 540152 425808 540204 425814
rect 540152 425750 540204 425756
rect 540164 419914 540192 425750
rect 540532 419914 540560 428606
rect 541164 427236 541216 427242
rect 541164 427178 541216 427184
rect 540980 423972 541032 423978
rect 540980 423914 541032 423920
rect 540992 419914 541020 423914
rect 541176 419914 541204 427178
rect 541348 420436 541400 420442
rect 541348 420378 541400 420384
rect 541360 420034 541388 420378
rect 541348 420028 541400 420034
rect 541348 419970 541400 419976
rect 541544 419914 541572 428742
rect 542360 425740 542412 425746
rect 542360 425682 542412 425688
rect 541900 423836 541952 423842
rect 541900 423778 541952 423784
rect 541624 420436 541676 420442
rect 541624 420378 541676 420384
rect 541636 420306 541664 420378
rect 541624 420300 541676 420306
rect 541624 420242 541676 420248
rect 541912 419914 541940 423778
rect 542372 419914 542400 425682
rect 542648 419914 542676 599558
rect 543016 425066 543044 700402
rect 543832 700392 543884 700398
rect 543832 700334 543884 700340
rect 543280 427168 543332 427174
rect 543280 427110 543332 427116
rect 543096 425128 543148 425134
rect 543096 425070 543148 425076
rect 543004 425060 543056 425066
rect 543004 425002 543056 425008
rect 542728 420640 542780 420646
rect 542728 420582 542780 420588
rect 542740 420306 542768 420582
rect 542728 420300 542780 420306
rect 542728 420242 542780 420248
rect 543108 419914 543136 425070
rect 543292 425054 543320 427110
rect 543740 425060 543792 425066
rect 543292 425026 543688 425054
rect 543660 419914 543688 425026
rect 543740 425002 543792 425008
rect 539888 419886 540086 419914
rect 540164 419886 540454 419914
rect 540532 419886 540822 419914
rect 540992 419886 541098 419914
rect 541176 419886 541466 419914
rect 541544 419886 541834 419914
rect 541912 419886 542202 419914
rect 542372 419886 542570 419914
rect 542648 419886 542938 419914
rect 543108 419886 543214 419914
rect 543598 419886 543688 419914
rect 543752 419914 543780 425002
rect 543844 423842 543872 700334
rect 543924 700324 543976 700330
rect 543924 700266 543976 700272
rect 543936 441614 543964 700266
rect 545304 670744 545356 670750
rect 545304 670686 545356 670692
rect 545212 656940 545264 656946
rect 545212 656882 545264 656888
rect 544384 618316 544436 618322
rect 544384 618258 544436 618264
rect 543936 441586 544332 441614
rect 544304 423858 544332 441586
rect 544396 423978 544424 618258
rect 545224 427814 545252 656882
rect 545316 441614 545344 670686
rect 554044 643136 554096 643142
rect 554044 643078 554096 643084
rect 546776 605872 546828 605878
rect 546776 605814 546828 605820
rect 546592 579692 546644 579698
rect 546592 579634 546644 579640
rect 545316 441586 545804 441614
rect 545224 427786 545436 427814
rect 544384 423972 544436 423978
rect 544384 423914 544436 423920
rect 543832 423836 543884 423842
rect 544304 423830 544424 423858
rect 543832 423778 543884 423784
rect 544014 422920 544070 422929
rect 544014 422855 544070 422864
rect 544028 419914 544056 422855
rect 544396 419914 544424 423830
rect 544752 423836 544804 423842
rect 544752 423778 544804 423784
rect 544764 419914 544792 423778
rect 545408 419914 545436 427786
rect 545776 419914 545804 441586
rect 546132 423904 546184 423910
rect 546132 423846 546184 423852
rect 546144 419914 546172 423846
rect 546604 423842 546632 579634
rect 546684 553444 546736 553450
rect 546684 553386 546736 553392
rect 546696 423910 546724 553386
rect 546788 441614 546816 605814
rect 548156 527196 548208 527202
rect 548156 527138 548208 527144
rect 547972 501016 548024 501022
rect 547972 500958 548024 500964
rect 546788 441586 546908 441614
rect 546684 423904 546736 423910
rect 546684 423846 546736 423852
rect 546592 423836 546644 423842
rect 546592 423778 546644 423784
rect 546684 420368 546736 420374
rect 546684 420310 546736 420316
rect 546592 420164 546644 420170
rect 546592 420106 546644 420112
rect 543752 419886 543950 419914
rect 544028 419886 544318 419914
rect 544396 419886 544686 419914
rect 544764 419886 544962 419914
rect 545408 419886 545698 419914
rect 545776 419886 546066 419914
rect 546144 419886 546434 419914
rect 546604 419830 546632 420106
rect 546696 419830 546724 420310
rect 546880 419914 546908 441586
rect 546960 423972 547012 423978
rect 546960 423914 547012 423920
rect 546818 419886 546908 419914
rect 546972 419914 547000 423914
rect 547512 423904 547564 423910
rect 547512 423846 547564 423852
rect 547144 423836 547196 423842
rect 547144 423778 547196 423784
rect 547156 419914 547184 423778
rect 547524 419914 547552 423846
rect 547984 423842 548012 500958
rect 548168 441614 548196 527138
rect 548168 441586 548288 441614
rect 548064 428528 548116 428534
rect 548064 428470 548116 428476
rect 547972 423836 548024 423842
rect 547972 423778 548024 423784
rect 547788 423156 547840 423162
rect 547788 423098 547840 423104
rect 547800 420374 547828 423098
rect 547972 420436 548024 420442
rect 547972 420378 548024 420384
rect 547788 420368 547840 420374
rect 547788 420310 547840 420316
rect 546972 419886 547078 419914
rect 547156 419886 547446 419914
rect 547524 419886 547814 419914
rect 547984 419898 548012 420378
rect 548076 419914 548104 428470
rect 548260 419914 548288 441586
rect 548892 428596 548944 428602
rect 548892 428538 548944 428544
rect 548616 423836 548668 423842
rect 548616 423778 548668 423784
rect 548524 422748 548576 422754
rect 548524 422690 548576 422696
rect 548536 421938 548564 422690
rect 548524 421932 548576 421938
rect 548524 421874 548576 421880
rect 548628 419914 548656 423778
rect 548904 419914 548932 428538
rect 549996 428460 550048 428466
rect 549996 428402 550048 428408
rect 549628 427100 549680 427106
rect 549628 427042 549680 427048
rect 549352 425196 549404 425202
rect 549352 425138 549404 425144
rect 549260 422884 549312 422890
rect 549260 422826 549312 422832
rect 549272 420442 549300 422826
rect 549260 420436 549312 420442
rect 549260 420378 549312 420384
rect 549364 419914 549392 425138
rect 549640 419914 549668 427042
rect 550008 419914 550036 428402
rect 554056 427514 554084 643078
rect 554044 427508 554096 427514
rect 554044 427450 554096 427456
rect 558932 424590 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580276 425950 580304 670647
rect 580354 564360 580410 564369
rect 580354 564295 580410 564304
rect 580264 425944 580316 425950
rect 580264 425886 580316 425892
rect 558920 424584 558972 424590
rect 558920 424526 558972 424532
rect 580368 424522 580396 564295
rect 580446 537840 580502 537849
rect 580446 537775 580502 537784
rect 580460 427446 580488 537775
rect 580538 511320 580594 511329
rect 580538 511255 580594 511264
rect 580448 427440 580500 427446
rect 580448 427382 580500 427388
rect 580356 424516 580408 424522
rect 580356 424458 580408 424464
rect 580552 424454 580580 511255
rect 580540 424448 580592 424454
rect 580540 424390 580592 424396
rect 556988 423768 557040 423774
rect 556988 423710 557040 423716
rect 550364 423564 550416 423570
rect 550364 423506 550416 423512
rect 550376 419914 550404 423506
rect 553584 423088 553636 423094
rect 551374 423056 551430 423065
rect 553584 423030 553636 423036
rect 551374 422991 551430 423000
rect 552204 423020 552256 423026
rect 551008 422952 551060 422958
rect 551008 422894 551060 422900
rect 550640 422340 550692 422346
rect 550640 422282 550692 422288
rect 550652 421705 550680 422282
rect 550638 421696 550694 421705
rect 550638 421631 550694 421640
rect 550640 421592 550692 421598
rect 550640 421534 550692 421540
rect 550652 419914 550680 421534
rect 551020 419914 551048 422894
rect 551388 419914 551416 422991
rect 552204 422962 552256 422968
rect 552110 420200 552166 420209
rect 552110 420135 552166 420144
rect 552124 419914 552152 420135
rect 547972 419892 548024 419898
rect 548076 419886 548182 419914
rect 548260 419886 548550 419914
rect 548628 419886 548826 419914
rect 548904 419886 549194 419914
rect 549364 419886 549562 419914
rect 549640 419886 549930 419914
rect 550008 419886 550298 419914
rect 550376 419886 550574 419914
rect 550652 419886 550942 419914
rect 551020 419886 551310 419914
rect 551388 419886 551678 419914
rect 552062 419886 552152 419914
rect 552216 419914 552244 422962
rect 552754 420336 552810 420345
rect 552754 420271 552810 420280
rect 552570 419928 552626 419937
rect 552216 419886 552414 419914
rect 552768 419914 552796 420271
rect 552626 419886 552690 419914
rect 552768 419886 553058 419914
rect 552570 419863 552626 419872
rect 547972 419834 548024 419840
rect 528142 419750 528416 419766
rect 529032 419750 529230 419778
rect 530626 419750 530808 419778
rect 534122 419750 534396 419778
rect 545212 419824 545264 419830
rect 546592 419824 546644 419830
rect 545264 419772 545330 419778
rect 545212 419766 545330 419772
rect 546592 419766 546644 419772
rect 546684 419824 546736 419830
rect 553596 419778 553624 423030
rect 556158 422784 556214 422793
rect 556158 422719 556214 422728
rect 554228 422544 554280 422550
rect 554228 422486 554280 422492
rect 554870 422512 554926 422521
rect 553858 421560 553914 421569
rect 553858 421495 553914 421504
rect 553676 420232 553728 420238
rect 553676 420174 553728 420180
rect 553688 419914 553716 420174
rect 553872 419914 553900 421495
rect 554240 419914 554268 422486
rect 554870 422447 554926 422456
rect 554884 419914 554912 422447
rect 555238 422376 555294 422385
rect 555238 422311 555294 422320
rect 555252 419914 555280 422311
rect 555700 419960 555752 419966
rect 553688 419886 553794 419914
rect 553872 419886 554162 419914
rect 554240 419886 554438 419914
rect 554884 419886 555174 419914
rect 555252 419886 555542 419914
rect 556172 419914 556200 422719
rect 556342 422648 556398 422657
rect 556342 422583 556398 422592
rect 556356 419914 556384 422583
rect 557000 419914 557028 423710
rect 557538 423192 557594 423201
rect 557538 423127 557594 423136
rect 557552 419914 557580 423127
rect 561036 422816 561088 422822
rect 561036 422758 561088 422764
rect 558368 422680 558420 422686
rect 558368 422622 558420 422628
rect 558092 422340 558144 422346
rect 558092 422282 558144 422288
rect 557814 420064 557870 420073
rect 557814 419999 557870 420008
rect 557828 419914 557856 419999
rect 558104 419914 558132 422282
rect 558380 419914 558408 422622
rect 560668 421864 560720 421870
rect 560668 421806 560720 421812
rect 560574 421288 560630 421297
rect 560574 421223 560630 421232
rect 560482 421152 560538 421161
rect 560482 421087 560538 421096
rect 560206 421016 560262 421025
rect 560206 420951 560262 420960
rect 559944 420022 560156 420050
rect 559194 419928 559250 419937
rect 555752 419908 555910 419914
rect 555700 419902 555910 419908
rect 555712 419886 555910 419902
rect 556172 419886 556278 419914
rect 556356 419886 556554 419914
rect 557000 419886 557290 419914
rect 557552 419886 557658 419914
rect 557828 419886 558026 419914
rect 558104 419886 558302 419914
rect 558380 419886 558670 419914
rect 559944 419914 559972 420022
rect 559250 419886 559406 419914
rect 559774 419886 559972 419914
rect 559194 419863 559250 419872
rect 546684 419766 546736 419772
rect 545224 419750 545330 419766
rect 553442 419750 553624 419778
rect 554596 419824 554648 419830
rect 556712 419824 556764 419830
rect 554648 419772 554806 419778
rect 554596 419766 554806 419772
rect 559288 419824 559340 419830
rect 556764 419772 556922 419778
rect 556712 419766 556922 419772
rect 554608 419750 554806 419766
rect 556724 419750 556922 419766
rect 559054 419772 559288 419778
rect 559054 419766 559340 419772
rect 559932 419824 559984 419830
rect 559932 419766 559984 419772
rect 560024 419824 560076 419830
rect 560024 419766 560076 419772
rect 559054 419750 559328 419766
rect 517518 419656 517574 419665
rect 517518 419591 517574 419600
rect 519820 419620 519872 419626
rect 517532 419558 517560 419591
rect 519820 419562 519872 419568
rect 514668 419552 514720 419558
rect 514668 419494 514720 419500
rect 517520 419552 517572 419558
rect 517520 419494 517572 419500
rect 447600 416900 447652 416906
rect 447600 416842 447652 416848
rect 447048 393372 447100 393378
rect 447048 393314 447100 393320
rect 446956 392012 447008 392018
rect 446956 391954 447008 391960
rect 446864 390584 446916 390590
rect 446864 390526 446916 390532
rect 446772 389224 446824 389230
rect 446772 389166 446824 389172
rect 446680 387932 446732 387938
rect 446680 387874 446732 387880
rect 446588 387864 446640 387870
rect 446588 387806 446640 387812
rect 446496 386436 446548 386442
rect 446496 386378 446548 386384
rect 446508 298110 446536 386378
rect 446496 298104 446548 298110
rect 446496 298046 446548 298052
rect 446600 297770 446628 387806
rect 446588 297764 446640 297770
rect 446588 297706 446640 297712
rect 446692 297702 446720 387874
rect 446784 297838 446812 389166
rect 446876 297906 446904 390526
rect 446968 297974 446996 391954
rect 446956 297968 447008 297974
rect 446956 297910 447008 297916
rect 446864 297900 446916 297906
rect 446864 297842 446916 297848
rect 446772 297832 446824 297838
rect 446772 297774 446824 297780
rect 446680 297696 446732 297702
rect 446680 297638 446732 297644
rect 447060 297634 447088 393314
rect 447612 365265 447640 416842
rect 447876 416832 447928 416838
rect 447876 416774 447928 416780
rect 447692 409896 447744 409902
rect 447692 409838 447744 409844
rect 447598 365256 447654 365265
rect 447598 365191 447654 365200
rect 447704 355473 447732 409838
rect 447784 404388 447836 404394
rect 447784 404330 447836 404336
rect 447690 355464 447746 355473
rect 447690 355399 447746 355408
rect 447796 345817 447824 404330
rect 447888 367169 447916 416774
rect 448980 415472 449032 415478
rect 448980 415414 449032 415420
rect 448152 392148 448204 392154
rect 448152 392090 448204 392096
rect 447968 392080 448020 392086
rect 447968 392022 448020 392028
rect 447874 367160 447930 367169
rect 447874 367095 447930 367104
rect 447874 366480 447930 366489
rect 447874 366415 447930 366424
rect 447782 345808 447838 345817
rect 447782 345743 447838 345752
rect 447782 302968 447838 302977
rect 447782 302903 447838 302912
rect 447048 297628 447100 297634
rect 447048 297570 447100 297576
rect 445668 200864 445720 200870
rect 445668 200806 445720 200812
rect 445484 200796 445536 200802
rect 445484 200738 445536 200744
rect 438124 200252 438176 200258
rect 438124 200194 438176 200200
rect 261576 167000 261628 167006
rect 261576 166942 261628 166948
rect 438136 86970 438164 200194
rect 438124 86964 438176 86970
rect 438124 86906 438176 86912
rect 447796 78810 447824 302903
rect 447888 301073 447916 366415
rect 447980 326233 448008 392022
rect 448060 390652 448112 390658
rect 448060 390594 448112 390600
rect 447966 326224 448022 326233
rect 447966 326159 448022 326168
rect 448072 322425 448100 390594
rect 448164 324329 448192 392090
rect 448244 389292 448296 389298
rect 448244 389234 448296 389240
rect 448150 324320 448206 324329
rect 448150 324255 448206 324264
rect 448058 322416 448114 322425
rect 448058 322351 448114 322360
rect 448256 320521 448284 389234
rect 448336 388000 448388 388006
rect 448336 387942 448388 387948
rect 448242 320512 448298 320521
rect 448242 320447 448298 320456
rect 448348 318481 448376 387942
rect 448428 386504 448480 386510
rect 448428 386446 448480 386452
rect 448334 318472 448390 318481
rect 448334 318407 448390 318416
rect 448440 316577 448468 386446
rect 448992 363225 449020 415414
rect 449072 414044 449124 414050
rect 449072 413986 449124 413992
rect 448978 363216 449034 363225
rect 448978 363151 449034 363160
rect 449084 361321 449112 413986
rect 450360 412684 450412 412690
rect 450360 412626 450412 412632
rect 450268 411324 450320 411330
rect 450268 411266 450320 411272
rect 450176 408536 450228 408542
rect 450176 408478 450228 408484
rect 449992 407244 450044 407250
rect 449992 407186 450044 407192
rect 449900 405748 449952 405754
rect 449900 405690 449952 405696
rect 449164 403028 449216 403034
rect 449164 402970 449216 402976
rect 449070 361312 449126 361321
rect 449070 361247 449126 361256
rect 449176 343777 449204 402970
rect 449348 401668 449400 401674
rect 449348 401610 449400 401616
rect 449256 400240 449308 400246
rect 449256 400182 449308 400188
rect 449162 343768 449218 343777
rect 449162 343703 449218 343712
rect 449268 339969 449296 400182
rect 449360 341873 449388 401610
rect 449532 400308 449584 400314
rect 449532 400250 449584 400256
rect 449440 397520 449492 397526
rect 449440 397462 449492 397468
rect 449346 341864 449402 341873
rect 449346 341799 449402 341808
rect 449254 339960 449310 339969
rect 449254 339895 449310 339904
rect 449452 334121 449480 397462
rect 449544 337929 449572 400250
rect 449624 398880 449676 398886
rect 449624 398822 449676 398828
rect 449530 337920 449586 337929
rect 449530 337855 449586 337864
rect 449636 336025 449664 398822
rect 449716 396092 449768 396098
rect 449716 396034 449768 396040
rect 449622 336016 449678 336025
rect 449622 335951 449678 335960
rect 449438 334112 449494 334121
rect 449438 334047 449494 334056
rect 449728 332081 449756 396034
rect 449808 394732 449860 394738
rect 449808 394674 449860 394680
rect 449714 332072 449770 332081
rect 449714 332007 449770 332016
rect 449820 330177 449848 394674
rect 449912 347857 449940 405690
rect 450004 350169 450032 407186
rect 450084 407176 450136 407182
rect 450084 407118 450136 407124
rect 450096 351937 450124 407118
rect 450188 354113 450216 408478
rect 450280 357649 450308 411266
rect 450372 359961 450400 412626
rect 450820 394800 450872 394806
rect 450820 394742 450872 394748
rect 450728 370524 450780 370530
rect 450728 370466 450780 370472
rect 450740 369617 450768 370466
rect 450726 369608 450782 369617
rect 450726 369543 450782 369552
rect 450358 359952 450414 359961
rect 450358 359887 450414 359896
rect 450266 357640 450322 357649
rect 450266 357575 450322 357584
rect 450174 354104 450230 354113
rect 450174 354039 450230 354048
rect 450082 351928 450138 351937
rect 450082 351863 450138 351872
rect 449990 350160 450046 350169
rect 449990 350095 450046 350104
rect 449898 347848 449954 347857
rect 449898 347783 449954 347792
rect 449806 330168 449862 330177
rect 449806 330103 449862 330112
rect 448426 316568 448482 316577
rect 448426 316503 448482 316512
rect 447874 301064 447930 301073
rect 447874 300999 447930 301008
rect 447784 78804 447836 78810
rect 447784 78746 447836 78752
rect 447888 78742 447916 300999
rect 450832 298042 450860 394742
rect 514022 385792 514078 385801
rect 514022 385727 514078 385736
rect 514036 385121 514064 385727
rect 514022 385112 514078 385121
rect 514022 385047 514078 385056
rect 509974 384704 510030 384713
rect 509974 384639 510030 384648
rect 509988 383761 510016 384639
rect 510158 384024 510214 384033
rect 510158 383959 510214 383968
rect 510172 383761 510200 383959
rect 509974 383752 510030 383761
rect 509974 383687 510030 383696
rect 510158 383752 510214 383761
rect 510158 383687 510214 383696
rect 514680 370598 514708 419494
rect 518162 419112 518218 419121
rect 518162 419047 518218 419056
rect 517610 417888 517666 417897
rect 517610 417823 517666 417832
rect 517520 416900 517572 416906
rect 517520 416842 517572 416848
rect 517532 416809 517560 416842
rect 517624 416838 517652 417823
rect 517612 416832 517664 416838
rect 517518 416800 517574 416809
rect 517612 416774 517664 416780
rect 517518 416735 517574 416744
rect 517518 415576 517574 415585
rect 517518 415511 517574 415520
rect 517532 415478 517560 415511
rect 517520 415472 517572 415478
rect 517520 415414 517572 415420
rect 517518 414352 517574 414361
rect 517518 414287 517574 414296
rect 517532 414050 517560 414287
rect 517520 414044 517572 414050
rect 517520 413986 517572 413992
rect 517518 413264 517574 413273
rect 517518 413199 517574 413208
rect 517532 412690 517560 413199
rect 517520 412684 517572 412690
rect 517520 412626 517572 412632
rect 517518 412040 517574 412049
rect 517518 411975 517574 411984
rect 517532 411330 517560 411975
rect 517794 411496 517850 411505
rect 517794 411431 517850 411440
rect 517520 411324 517572 411330
rect 517520 411266 517572 411272
rect 517518 410816 517574 410825
rect 517518 410751 517574 410760
rect 517532 409902 517560 410751
rect 517520 409896 517572 409902
rect 517520 409838 517572 409844
rect 517518 409728 517574 409737
rect 517518 409663 517574 409672
rect 517532 408542 517560 409663
rect 517520 408536 517572 408542
rect 517520 408478 517572 408484
rect 517610 408504 517666 408513
rect 517610 408439 517666 408448
rect 517518 407280 517574 407289
rect 517518 407215 517520 407224
rect 517572 407215 517574 407224
rect 517520 407186 517572 407192
rect 517624 407182 517652 408439
rect 517612 407176 517664 407182
rect 517612 407118 517664 407124
rect 517518 406192 517574 406201
rect 517518 406127 517574 406136
rect 517532 405754 517560 406127
rect 517520 405748 517572 405754
rect 517520 405690 517572 405696
rect 517518 404968 517574 404977
rect 517518 404903 517574 404912
rect 517532 404394 517560 404903
rect 517520 404388 517572 404394
rect 517520 404330 517572 404336
rect 517808 404274 517836 411431
rect 517886 407960 517942 407969
rect 517886 407895 517942 407904
rect 517532 404246 517836 404274
rect 517532 370870 517560 404246
rect 517900 404138 517928 407895
rect 517624 404110 517928 404138
rect 517624 379914 517652 404110
rect 517702 403744 517758 403753
rect 517702 403679 517758 403688
rect 517716 403034 517744 403679
rect 517704 403028 517756 403034
rect 517704 402970 517756 402976
rect 517702 402656 517758 402665
rect 517702 402591 517758 402600
rect 517716 401674 517744 402591
rect 517704 401668 517756 401674
rect 517704 401610 517756 401616
rect 517794 401432 517850 401441
rect 517794 401367 517850 401376
rect 517702 400344 517758 400353
rect 517702 400279 517704 400288
rect 517756 400279 517758 400288
rect 517704 400250 517756 400256
rect 517808 400246 517836 401367
rect 517796 400240 517848 400246
rect 517796 400182 517848 400188
rect 517702 399120 517758 399129
rect 517702 399055 517758 399064
rect 517716 398886 517744 399055
rect 517704 398880 517756 398886
rect 517704 398822 517756 398828
rect 517702 397896 517758 397905
rect 517702 397831 517758 397840
rect 517716 397526 517744 397831
rect 517704 397520 517756 397526
rect 517704 397462 517756 397468
rect 517702 396808 517758 396817
rect 517702 396743 517758 396752
rect 517716 396098 517744 396743
rect 517886 396128 517942 396137
rect 517704 396092 517756 396098
rect 517886 396063 517942 396072
rect 517704 396034 517756 396040
rect 517794 395584 517850 395593
rect 517794 395519 517850 395528
rect 517702 395040 517758 395049
rect 517702 394975 517758 394984
rect 517716 394806 517744 394975
rect 517704 394800 517756 394806
rect 517704 394742 517756 394748
rect 517808 394738 517836 395519
rect 517796 394732 517848 394738
rect 517796 394674 517848 394680
rect 517900 394618 517928 396063
rect 517808 394590 517928 394618
rect 517702 393816 517758 393825
rect 517702 393751 517758 393760
rect 517716 393378 517744 393751
rect 517704 393372 517756 393378
rect 517704 393314 517756 393320
rect 517704 392148 517756 392154
rect 517704 392090 517756 392096
rect 517716 392057 517744 392090
rect 517702 392048 517758 392057
rect 517702 391983 517758 391992
rect 517702 390824 517758 390833
rect 517702 390759 517758 390768
rect 517716 390658 517744 390759
rect 517704 390652 517756 390658
rect 517704 390594 517756 390600
rect 517702 389736 517758 389745
rect 517702 389671 517758 389680
rect 517716 389298 517744 389671
rect 517704 389292 517756 389298
rect 517704 389234 517756 389240
rect 517702 387968 517758 387977
rect 517702 387903 517704 387912
rect 517756 387903 517758 387912
rect 517704 387874 517756 387880
rect 517702 386744 517758 386753
rect 517702 386679 517758 386688
rect 517716 386442 517744 386679
rect 517704 386436 517756 386442
rect 517704 386378 517756 386384
rect 517612 379908 517664 379914
rect 517612 379850 517664 379856
rect 517808 379001 517836 394590
rect 517886 393272 517942 393281
rect 517886 393207 517942 393216
rect 517900 392086 517928 393207
rect 517978 392592 518034 392601
rect 517978 392527 518034 392536
rect 517888 392080 517940 392086
rect 517888 392022 517940 392028
rect 517992 392018 518020 392527
rect 517980 392012 518032 392018
rect 517980 391954 518032 391960
rect 517886 391504 517942 391513
rect 517886 391439 517942 391448
rect 517900 390590 517928 391439
rect 517888 390584 517940 390590
rect 517888 390526 517940 390532
rect 517886 390280 517942 390289
rect 517886 390215 517942 390224
rect 517900 389230 517928 390215
rect 517888 389224 517940 389230
rect 517888 389166 517940 389172
rect 517978 389056 518034 389065
rect 517978 388991 518034 389000
rect 517886 388512 517942 388521
rect 517886 388447 517942 388456
rect 517900 388006 517928 388447
rect 517888 388000 517940 388006
rect 517888 387942 517940 387948
rect 517992 387870 518020 388991
rect 517980 387864 518032 387870
rect 517980 387806 518032 387812
rect 517886 387288 517942 387297
rect 517886 387223 517942 387232
rect 517900 386510 517928 387223
rect 517888 386504 517940 386510
rect 517888 386446 517940 386452
rect 518070 380896 518126 380905
rect 518070 380831 518126 380840
rect 517794 378992 517850 379001
rect 517794 378927 517850 378936
rect 518084 372065 518112 380831
rect 518070 372056 518126 372065
rect 518070 371991 518126 372000
rect 517520 370864 517572 370870
rect 517520 370806 517572 370812
rect 514668 370592 514720 370598
rect 514668 370534 514720 370540
rect 518176 370530 518204 419047
rect 519832 419014 519860 419562
rect 519910 419384 519966 419393
rect 519966 419342 520122 419370
rect 519910 419319 519966 419328
rect 519820 419008 519872 419014
rect 519820 418950 519872 418956
rect 518806 417344 518862 417353
rect 518806 417279 518862 417288
rect 518714 416120 518770 416129
rect 518714 416055 518770 416064
rect 518622 415032 518678 415041
rect 518622 414967 518678 414976
rect 518530 413808 518586 413817
rect 518530 413743 518586 413752
rect 518346 412584 518402 412593
rect 518346 412519 518402 412528
rect 518254 410272 518310 410281
rect 518254 410207 518310 410216
rect 518268 370802 518296 410207
rect 518256 370796 518308 370802
rect 518256 370738 518308 370744
rect 518360 370705 518388 412519
rect 518544 370977 518572 413743
rect 518530 370968 518586 370977
rect 518530 370903 518586 370912
rect 518346 370696 518402 370705
rect 518346 370631 518402 370640
rect 518636 370530 518664 414967
rect 518728 370734 518756 416055
rect 518716 370728 518768 370734
rect 518716 370670 518768 370676
rect 518820 370666 518848 417279
rect 518898 409048 518954 409057
rect 518898 408983 518954 408992
rect 518912 370938 518940 408983
rect 518990 406736 519046 406745
rect 518990 406671 519046 406680
rect 519004 379030 519032 406671
rect 519266 405512 519322 405521
rect 519266 405447 519322 405456
rect 519082 404424 519138 404433
rect 519082 404359 519138 404368
rect 519096 379098 519124 404359
rect 519174 403200 519230 403209
rect 519174 403135 519230 403144
rect 519084 379092 519136 379098
rect 519084 379034 519136 379040
rect 518992 379024 519044 379030
rect 518992 378966 519044 378972
rect 519188 378894 519216 403135
rect 519176 378888 519228 378894
rect 519176 378830 519228 378836
rect 519280 378826 519308 405447
rect 519358 401976 519414 401985
rect 519358 401911 519414 401920
rect 519372 379166 519400 401911
rect 519450 400888 519506 400897
rect 519450 400823 519506 400832
rect 519360 379160 519412 379166
rect 519360 379102 519412 379108
rect 519464 378962 519492 400823
rect 519542 399664 519598 399673
rect 519542 399599 519598 399608
rect 519556 379137 519584 399599
rect 519726 398576 519782 398585
rect 519726 398511 519782 398520
rect 519542 379128 519598 379137
rect 519542 379063 519598 379072
rect 519452 378956 519504 378962
rect 519452 378898 519504 378904
rect 519740 378865 519768 398511
rect 519726 378856 519782 378865
rect 519268 378820 519320 378826
rect 519726 378791 519782 378800
rect 519268 378762 519320 378768
rect 520108 374678 520136 380052
rect 520384 377466 520412 380037
rect 520372 377460 520424 377466
rect 520372 377402 520424 377408
rect 520660 374746 520688 380037
rect 520648 374740 520700 374746
rect 520648 374682 520700 374688
rect 520096 374672 520148 374678
rect 520096 374614 520148 374620
rect 521028 371890 521056 380037
rect 521304 377738 521332 380037
rect 521580 378078 521608 380037
rect 521568 378072 521620 378078
rect 521568 378014 521620 378020
rect 521292 377732 521344 377738
rect 521292 377674 521344 377680
rect 521016 371884 521068 371890
rect 521016 371826 521068 371832
rect 521948 371006 521976 380037
rect 522224 371074 522252 380037
rect 522500 371142 522528 380037
rect 522868 371210 522896 380037
rect 523040 378072 523092 378078
rect 523040 378014 523092 378020
rect 523052 376038 523080 378014
rect 523144 376106 523172 380037
rect 523420 377602 523448 380037
rect 523408 377596 523460 377602
rect 523408 377538 523460 377544
rect 523132 376100 523184 376106
rect 523132 376042 523184 376048
rect 523040 376032 523092 376038
rect 523040 375974 523092 375980
rect 523788 374814 523816 380037
rect 524064 377534 524092 380037
rect 524340 377670 524368 380037
rect 524328 377664 524380 377670
rect 524328 377606 524380 377612
rect 524052 377528 524104 377534
rect 524052 377470 524104 377476
rect 524708 376174 524736 380037
rect 550640 379908 550692 379914
rect 550640 379850 550692 379856
rect 549628 379160 549680 379166
rect 549628 379102 549680 379108
rect 533344 377732 533396 377738
rect 533344 377674 533396 377680
rect 524696 376168 524748 376174
rect 524696 376110 524748 376116
rect 523776 374808 523828 374814
rect 523776 374750 523828 374756
rect 533356 371958 533384 377674
rect 549260 377460 549312 377466
rect 549260 377402 549312 377408
rect 533344 371952 533396 371958
rect 533344 371894 533396 371900
rect 522856 371204 522908 371210
rect 522856 371146 522908 371152
rect 522488 371136 522540 371142
rect 522488 371078 522540 371084
rect 522212 371068 522264 371074
rect 522212 371010 522264 371016
rect 521936 371000 521988 371006
rect 521936 370942 521988 370948
rect 518900 370932 518952 370938
rect 518900 370874 518952 370880
rect 518808 370660 518860 370666
rect 518808 370602 518860 370608
rect 518164 370524 518216 370530
rect 518164 370466 518216 370472
rect 518624 370524 518676 370530
rect 518624 370466 518676 370472
rect 549272 307170 549300 377402
rect 549352 371884 549404 371890
rect 549352 371826 549404 371832
rect 549364 315761 549392 371826
rect 549536 370932 549588 370938
rect 549536 370874 549588 370880
rect 549444 370864 549496 370870
rect 549444 370806 549496 370812
rect 549350 315752 549406 315761
rect 549350 315687 549406 315696
rect 549350 307184 549406 307193
rect 549272 307142 549350 307170
rect 549350 307119 549406 307128
rect 548366 300070 548656 300098
rect 451476 299577 451504 300037
rect 454540 299826 454568 300016
rect 457668 299826 457696 300016
rect 460796 299826 460824 300016
rect 454512 299798 454568 299826
rect 457640 299798 457696 299826
rect 460768 299798 460824 299826
rect 451462 299568 451518 299577
rect 451462 299503 451518 299512
rect 450820 298036 450872 298042
rect 450820 297978 450872 297984
rect 454512 297945 454540 299798
rect 454498 297936 454554 297945
rect 454498 297871 454554 297880
rect 457640 297809 457668 299798
rect 460768 298110 460796 299798
rect 463924 299792 463952 300016
rect 467052 299792 467080 300016
rect 470180 299792 470208 300016
rect 473308 299792 473336 300016
rect 476436 299792 476464 300016
rect 479564 299792 479592 300016
rect 482692 299826 482720 300016
rect 485820 299826 485848 300016
rect 488948 299826 488976 300016
rect 492076 299826 492104 300016
rect 495204 299826 495232 300016
rect 498332 299826 498360 300016
rect 501460 299826 501488 300016
rect 504588 299826 504616 300016
rect 507716 299826 507744 300016
rect 510844 299826 510872 300016
rect 513972 299826 514000 300016
rect 517100 299826 517128 300016
rect 520228 299826 520256 300016
rect 523356 299826 523384 300016
rect 526484 299826 526512 300016
rect 529612 299826 529640 300016
rect 532740 299826 532768 300016
rect 535868 299826 535896 300016
rect 538996 299826 539024 300016
rect 542124 299826 542152 300016
rect 545252 299826 545280 300016
rect 463896 299764 463952 299792
rect 467024 299764 467080 299792
rect 470152 299764 470208 299792
rect 473280 299764 473336 299792
rect 476408 299764 476464 299792
rect 479536 299764 479592 299792
rect 482664 299798 482720 299826
rect 485792 299798 485848 299826
rect 488920 299798 488976 299826
rect 492048 299798 492104 299826
rect 495176 299798 495232 299826
rect 498304 299798 498360 299826
rect 501432 299798 501488 299826
rect 504560 299798 504616 299826
rect 507688 299798 507744 299826
rect 510816 299798 510872 299826
rect 513944 299798 514000 299826
rect 517072 299798 517128 299826
rect 520200 299798 520256 299826
rect 523328 299798 523384 299826
rect 526456 299798 526512 299826
rect 529584 299798 529640 299826
rect 532712 299798 532768 299826
rect 535840 299798 535896 299826
rect 538968 299798 539024 299826
rect 542096 299798 542152 299826
rect 545224 299798 545280 299826
rect 460756 298104 460808 298110
rect 460756 298046 460808 298052
rect 457626 297800 457682 297809
rect 457626 297735 457682 297744
rect 463896 297702 463924 299764
rect 467024 297770 467052 299764
rect 470152 297838 470180 299764
rect 473280 297906 473308 299764
rect 476408 297974 476436 299764
rect 476396 297968 476448 297974
rect 476396 297910 476448 297916
rect 473268 297900 473320 297906
rect 473268 297842 473320 297848
rect 470140 297832 470192 297838
rect 470140 297774 470192 297780
rect 467012 297764 467064 297770
rect 467012 297706 467064 297712
rect 463884 297696 463936 297702
rect 463884 297638 463936 297644
rect 479536 297634 479564 299764
rect 482664 298042 482692 299798
rect 482652 298036 482704 298042
rect 482652 297978 482704 297984
rect 479524 297628 479576 297634
rect 479524 297570 479576 297576
rect 485792 297265 485820 299798
rect 488920 297945 488948 299798
rect 488906 297936 488962 297945
rect 488906 297871 488962 297880
rect 492048 297809 492076 299798
rect 492034 297800 492090 297809
rect 492034 297735 492090 297744
rect 495176 297673 495204 299798
rect 495162 297664 495218 297673
rect 495162 297599 495218 297608
rect 498304 297498 498332 299798
rect 498292 297492 498344 297498
rect 498292 297434 498344 297440
rect 501432 297430 501460 299798
rect 501420 297424 501472 297430
rect 501420 297366 501472 297372
rect 504560 297362 504588 299798
rect 504548 297356 504600 297362
rect 504548 297298 504600 297304
rect 507688 297294 507716 299798
rect 510816 297838 510844 299798
rect 510804 297832 510856 297838
rect 510804 297774 510856 297780
rect 513944 297770 513972 299798
rect 513932 297764 513984 297770
rect 513932 297706 513984 297712
rect 517072 297702 517100 299798
rect 517060 297696 517112 297702
rect 517060 297638 517112 297644
rect 520200 297634 520228 299798
rect 520188 297628 520240 297634
rect 520188 297570 520240 297576
rect 523328 297566 523356 299798
rect 523316 297560 523368 297566
rect 523316 297502 523368 297508
rect 507676 297288 507728 297294
rect 485778 297256 485834 297265
rect 507676 297230 507728 297236
rect 526456 297226 526484 299798
rect 529584 297401 529612 299798
rect 532712 297537 532740 299798
rect 535840 298042 535868 299798
rect 535828 298036 535880 298042
rect 535828 297978 535880 297984
rect 538968 297974 538996 299798
rect 538956 297968 539008 297974
rect 538956 297910 539008 297916
rect 542096 297906 542124 299798
rect 545224 298110 545252 299798
rect 545212 298104 545264 298110
rect 548628 298081 548656 300070
rect 545212 298046 545264 298052
rect 548614 298072 548670 298081
rect 548614 298007 548670 298016
rect 542084 297900 542136 297906
rect 542084 297842 542136 297848
rect 532698 297528 532754 297537
rect 532698 297463 532754 297472
rect 529570 297392 529626 297401
rect 529570 297327 529626 297336
rect 549456 297226 549484 370806
rect 549548 297634 549576 370874
rect 549536 297628 549588 297634
rect 549536 297570 549588 297576
rect 549640 297430 549668 379102
rect 549720 379092 549772 379098
rect 549720 379034 549772 379040
rect 549628 297424 549680 297430
rect 549628 297366 549680 297372
rect 549732 297294 549760 379034
rect 549812 379024 549864 379030
rect 549812 378966 549864 378972
rect 549824 297770 549852 378966
rect 549904 377664 549956 377670
rect 549904 377606 549956 377612
rect 549916 363905 549944 377606
rect 549996 377596 550048 377602
rect 549996 377538 550048 377544
rect 549902 363896 549958 363905
rect 549902 363831 549958 363840
rect 549904 352572 549956 352578
rect 549904 352514 549956 352520
rect 549812 297764 549864 297770
rect 549812 297706 549864 297712
rect 549720 297288 549772 297294
rect 549720 297230 549772 297236
rect 485778 297191 485834 297200
rect 526444 297220 526496 297226
rect 526444 297162 526496 297168
rect 549444 297220 549496 297226
rect 549444 297162 549496 297168
rect 549916 202162 549944 352514
rect 550008 350418 550036 377538
rect 550088 376168 550140 376174
rect 550088 376110 550140 376116
rect 550100 367849 550128 376110
rect 550086 367840 550142 367849
rect 550086 367775 550142 367784
rect 550086 350432 550142 350441
rect 550008 350390 550086 350418
rect 550086 350367 550142 350376
rect 550652 297702 550680 379850
rect 550732 378956 550784 378962
rect 550732 378898 550784 378904
rect 550640 297696 550692 297702
rect 550640 297638 550692 297644
rect 550744 297498 550772 378898
rect 550824 378888 550876 378894
rect 550824 378830 550876 378836
rect 550732 297492 550784 297498
rect 550732 297434 550784 297440
rect 550836 297362 550864 378830
rect 550916 378820 550968 378826
rect 550916 378762 550968 378768
rect 550928 297838 550956 378762
rect 551468 377528 551520 377534
rect 551468 377470 551520 377476
rect 551284 376100 551336 376106
rect 551284 376042 551336 376048
rect 551192 374740 551244 374746
rect 551192 374682 551244 374688
rect 551100 374672 551152 374678
rect 551100 374614 551152 374620
rect 551008 370796 551060 370802
rect 551008 370738 551060 370744
rect 550916 297832 550968 297838
rect 550916 297774 550968 297780
rect 551020 297566 551048 370738
rect 551112 302297 551140 374614
rect 551204 311001 551232 374682
rect 551296 345953 551324 376042
rect 551376 374808 551428 374814
rect 551376 374750 551428 374756
rect 551388 354793 551416 374750
rect 551480 359145 551508 377470
rect 552112 376032 552164 376038
rect 552112 375974 552164 375980
rect 552020 371952 552072 371958
rect 552020 371894 552072 371900
rect 551466 359136 551522 359145
rect 551466 359071 551522 359080
rect 551374 354784 551430 354793
rect 551374 354719 551430 354728
rect 551282 345944 551338 345953
rect 551282 345879 551338 345888
rect 552032 319705 552060 371894
rect 552124 324057 552152 375974
rect 552480 371204 552532 371210
rect 552480 371146 552532 371152
rect 552388 371136 552440 371142
rect 552388 371078 552440 371084
rect 552296 371068 552348 371074
rect 552296 371010 552348 371016
rect 552204 371000 552256 371006
rect 552204 370942 552256 370948
rect 552216 328545 552244 370942
rect 552308 332897 552336 371010
rect 552400 337249 552428 371078
rect 552492 341601 552520 371146
rect 553584 370728 553636 370734
rect 553584 370670 553636 370676
rect 553398 370560 553454 370569
rect 553398 370495 553454 370504
rect 553492 370524 553544 370530
rect 552478 341592 552534 341601
rect 552478 341527 552534 341536
rect 552386 337240 552442 337249
rect 552386 337175 552442 337184
rect 552294 332888 552350 332897
rect 552294 332823 552350 332832
rect 552202 328536 552258 328545
rect 552202 328471 552258 328480
rect 552110 324048 552166 324057
rect 552110 323983 552166 323992
rect 552018 319696 552074 319705
rect 552018 319631 552074 319640
rect 551190 310992 551246 311001
rect 551190 310927 551246 310936
rect 551098 302288 551154 302297
rect 551098 302223 551154 302232
rect 553412 298110 553440 370495
rect 553492 370466 553544 370472
rect 553400 298104 553452 298110
rect 553400 298046 553452 298052
rect 553504 298042 553532 370466
rect 553492 298036 553544 298042
rect 553492 297978 553544 297984
rect 553596 297974 553624 370670
rect 553676 370660 553728 370666
rect 553676 370602 553728 370608
rect 553584 297968 553636 297974
rect 553584 297910 553636 297916
rect 553688 297906 553716 370602
rect 553768 370592 553820 370598
rect 553768 370534 553820 370540
rect 553780 298081 553808 370534
rect 553766 298072 553822 298081
rect 553766 298007 553822 298016
rect 553676 297900 553728 297906
rect 553676 297842 553728 297848
rect 551008 297560 551060 297566
rect 551008 297502 551060 297508
rect 550824 297356 550876 297362
rect 550824 297298 550876 297304
rect 559944 202230 559972 419766
rect 559932 202224 559984 202230
rect 559932 202166 559984 202172
rect 549904 202156 549956 202162
rect 549904 202098 549956 202104
rect 560036 126954 560064 419766
rect 560024 126948 560076 126954
rect 560024 126890 560076 126896
rect 447876 78736 447928 78742
rect 447876 78678 447928 78684
rect 289084 78260 289136 78266
rect 289084 78202 289136 78208
rect 287060 75472 287112 75478
rect 287060 75414 287112 75420
rect 284300 74112 284352 74118
rect 284300 74054 284352 74060
rect 280160 72752 280212 72758
rect 280160 72694 280212 72700
rect 276020 71324 276072 71330
rect 276020 71266 276072 71272
rect 273260 69964 273312 69970
rect 273260 69906 273312 69912
rect 269120 68604 269172 68610
rect 269120 68546 269172 68552
rect 266360 67176 266412 67182
rect 266360 67118 266412 67124
rect 262220 65816 262272 65822
rect 262220 65758 262272 65764
rect 261484 46912 261536 46918
rect 261484 46854 261536 46860
rect 262232 16574 262260 65758
rect 264980 52012 265032 52018
rect 264980 51954 265032 51960
rect 263600 27192 263652 27198
rect 263600 27134 263652 27140
rect 263612 16574 263640 27134
rect 259656 16546 260696 16574
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 259472 3454 259592 3482
rect 259472 480 259500 3454
rect 260668 480 260696 16546
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264164 480 264192 16546
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 51954
rect 266372 16574 266400 67118
rect 267740 53440 267792 53446
rect 267740 53382 267792 53388
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267752 3602 267780 53382
rect 267832 28620 267884 28626
rect 267832 28562 267884 28568
rect 267740 3596 267792 3602
rect 267740 3538 267792 3544
rect 267844 3482 267872 28562
rect 269132 16574 269160 68546
rect 271880 53372 271932 53378
rect 271880 53314 271932 53320
rect 270500 41064 270552 41070
rect 270500 41006 270552 41012
rect 270512 16574 270540 41006
rect 271892 16574 271920 53314
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 268476 3596 268528 3602
rect 268476 3538 268528 3544
rect 267752 3454 267872 3482
rect 267752 480 267780 3454
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268488 354 268516 3538
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268488 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 69906
rect 274640 28552 274692 28558
rect 274640 28494 274692 28500
rect 274652 16574 274680 28494
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 276032 3602 276060 71266
rect 278780 56228 278832 56234
rect 278780 56170 278832 56176
rect 276112 54868 276164 54874
rect 276112 54810 276164 54816
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 276124 3482 276152 54810
rect 277400 29980 277452 29986
rect 277400 29922 277452 29928
rect 277412 16574 277440 29922
rect 278792 16574 278820 56170
rect 280172 16574 280200 72694
rect 282920 56160 282972 56166
rect 282920 56102 282972 56108
rect 281540 45144 281592 45150
rect 281540 45086 281592 45092
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 276756 3596 276808 3602
rect 276756 3538 276808 3544
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 3538
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 45086
rect 282932 16574 282960 56102
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 480 284340 74054
rect 285680 57588 285732 57594
rect 285680 57530 285732 57536
rect 284392 40996 284444 41002
rect 284392 40938 284444 40944
rect 284404 16574 284432 40938
rect 285692 16574 285720 57530
rect 287072 16574 287100 75414
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289096 6254 289124 78202
rect 418804 78192 418856 78198
rect 418804 78134 418856 78140
rect 407764 78056 407816 78062
rect 407764 77998 407816 78004
rect 291200 76832 291252 76838
rect 291200 76774 291252 76780
rect 289820 57520 289872 57526
rect 289820 57462 289872 57468
rect 288992 6248 289044 6254
rect 288992 6190 289044 6196
rect 289084 6248 289136 6254
rect 289084 6190 289136 6196
rect 289004 480 289032 6190
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 57462
rect 291212 16574 291240 76774
rect 374000 75404 374052 75410
rect 374000 75346 374052 75352
rect 357440 67108 357492 67114
rect 357440 67050 357492 67056
rect 346400 65748 346452 65754
rect 346400 65690 346452 65696
rect 335360 64388 335412 64394
rect 335360 64330 335412 64336
rect 293960 63096 294012 63102
rect 293960 63038 294012 63044
rect 292580 59016 292632 59022
rect 292580 58958 292632 58964
rect 292592 16574 292620 58958
rect 293972 16574 294000 63038
rect 324320 63028 324372 63034
rect 324320 62970 324372 62976
rect 314660 61668 314712 61674
rect 314660 61610 314712 61616
rect 303620 60308 303672 60314
rect 303620 60250 303672 60256
rect 296720 58948 296772 58954
rect 296720 58890 296772 58896
rect 295340 42356 295392 42362
rect 295340 42298 295392 42304
rect 295352 16574 295380 42298
rect 296732 16574 296760 58890
rect 298100 51944 298152 51950
rect 298100 51886 298152 51892
rect 291212 16546 291424 16574
rect 292592 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 291396 480 291424 16546
rect 292580 6452 292632 6458
rect 292580 6394 292632 6400
rect 292592 480 292620 6394
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 51886
rect 302240 29912 302292 29918
rect 302240 29854 302292 29860
rect 300860 20256 300912 20262
rect 300860 20198 300912 20204
rect 300872 16574 300900 20198
rect 302252 16574 302280 29854
rect 303632 16574 303660 60250
rect 307760 60240 307812 60246
rect 307760 60182 307812 60188
rect 306380 31340 306432 31346
rect 306380 31282 306432 31288
rect 305000 20188 305052 20194
rect 305000 20130 305052 20136
rect 305012 16574 305040 20130
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299480 13388 299532 13394
rect 299480 13330 299532 13336
rect 299492 2786 299520 13330
rect 299664 6384 299716 6390
rect 299664 6326 299716 6332
rect 299480 2780 299532 2786
rect 299480 2722 299532 2728
rect 299676 480 299704 6326
rect 300768 2780 300820 2786
rect 300768 2722 300820 2728
rect 300780 480 300808 2722
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 31282
rect 307772 3482 307800 60182
rect 310520 60172 310572 60178
rect 310520 60114 310572 60120
rect 309140 31272 309192 31278
rect 309140 31214 309192 31220
rect 307852 20120 307904 20126
rect 307852 20062 307904 20068
rect 307864 3602 307892 20062
rect 309152 16574 309180 31214
rect 310532 16574 310560 60114
rect 313280 31204 313332 31210
rect 313280 31146 313332 31152
rect 311900 20052 311952 20058
rect 311900 19994 311952 20000
rect 311912 16574 311940 19994
rect 313292 16574 313320 31146
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 307852 3596 307904 3602
rect 307852 3538 307904 3544
rect 309048 3596 309100 3602
rect 309048 3538 309100 3544
rect 307772 3454 307984 3482
rect 307956 480 307984 3454
rect 309060 480 309088 3538
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311452 480 311480 16546
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 61610
rect 317420 61600 317472 61606
rect 317420 61542 317472 61548
rect 316040 32700 316092 32706
rect 316040 32642 316092 32648
rect 316052 3602 316080 32642
rect 317432 16574 317460 61542
rect 321560 61532 321612 61538
rect 321560 61474 321612 61480
rect 320180 32632 320232 32638
rect 320180 32574 320232 32580
rect 318800 21684 318852 21690
rect 318800 21626 318852 21632
rect 318812 16574 318840 21626
rect 320192 16574 320220 32574
rect 321572 16574 321600 61474
rect 322940 18896 322992 18902
rect 322940 18838 322992 18844
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316224 12028 316276 12034
rect 316224 11970 316276 11976
rect 316040 3596 316092 3602
rect 316040 3538 316092 3544
rect 316236 480 316264 11970
rect 317328 3596 317380 3602
rect 317328 3538 317380 3544
rect 317340 480 317368 3538
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 18838
rect 324332 3602 324360 62970
rect 328460 62960 328512 62966
rect 328460 62902 328512 62908
rect 327080 34060 327132 34066
rect 327080 34002 327132 34008
rect 324412 32564 324464 32570
rect 324412 32506 324464 32512
rect 324320 3596 324372 3602
rect 324320 3538 324372 3544
rect 324424 480 324452 32506
rect 325700 17536 325752 17542
rect 325700 17478 325752 17484
rect 325712 16574 325740 17478
rect 327092 16574 327120 34002
rect 328472 16574 328500 62902
rect 332600 62892 332652 62898
rect 332600 62834 332652 62840
rect 331220 33992 331272 33998
rect 331220 33934 331272 33940
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 325608 3596 325660 3602
rect 325608 3538 325660 3544
rect 325620 480 325648 3538
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330392 5092 330444 5098
rect 330392 5034 330444 5040
rect 330404 480 330432 5034
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 33934
rect 332612 3482 332640 62834
rect 333980 33924 334032 33930
rect 333980 33866 334032 33872
rect 332692 21616 332744 21622
rect 332692 21558 332744 21564
rect 332704 3602 332732 21558
rect 333992 16574 334020 33866
rect 335372 16574 335400 64330
rect 339500 64320 339552 64326
rect 339500 64262 339552 64268
rect 338120 35420 338172 35426
rect 338120 35362 338172 35368
rect 336740 21548 336792 21554
rect 336740 21490 336792 21496
rect 336752 16574 336780 21490
rect 338132 16574 338160 35362
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 332692 3596 332744 3602
rect 332692 3538 332744 3544
rect 333888 3596 333940 3602
rect 333888 3538 333940 3544
rect 332612 3454 332732 3482
rect 332704 480 332732 3454
rect 333900 480 333928 3538
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336292 480 336320 16546
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 64262
rect 342260 64252 342312 64258
rect 342260 64194 342312 64200
rect 340880 35488 340932 35494
rect 340880 35430 340932 35436
rect 340892 2378 340920 35430
rect 340972 21480 341024 21486
rect 340972 21422 341024 21428
rect 340880 2372 340932 2378
rect 340880 2314 340932 2320
rect 340984 480 341012 21422
rect 342272 16574 342300 64194
rect 345020 36848 345072 36854
rect 345020 36790 345072 36796
rect 343640 25764 343692 25770
rect 343640 25706 343692 25712
rect 343652 16574 343680 25706
rect 345032 16574 345060 36790
rect 346412 16574 346440 65690
rect 349160 65680 349212 65686
rect 349160 65622 349212 65628
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 342168 2372 342220 2378
rect 342168 2314 342220 2320
rect 342180 480 342208 2314
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348056 16176 348108 16182
rect 348056 16118 348108 16124
rect 348068 480 348096 16118
rect 349172 2378 349200 65622
rect 353300 65612 353352 65618
rect 353300 65554 353352 65560
rect 350540 28484 350592 28490
rect 350540 28426 350592 28432
rect 350552 16574 350580 28426
rect 353312 16574 353340 65554
rect 354680 49224 354732 49230
rect 354680 49166 354732 49172
rect 354692 16574 354720 49166
rect 356060 45076 356112 45082
rect 356060 45018 356112 45024
rect 356072 16574 356100 45018
rect 350552 16546 351224 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 349252 7880 349304 7886
rect 349252 7822 349304 7828
rect 349160 2372 349212 2378
rect 349160 2314 349212 2320
rect 349264 480 349292 7822
rect 350448 2372 350500 2378
rect 350448 2314 350500 2320
rect 350460 480 350488 2314
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352840 7812 352892 7818
rect 352840 7754 352892 7760
rect 352852 480 352880 7754
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357452 3482 357480 67050
rect 371240 67040 371292 67046
rect 371240 66982 371292 66988
rect 368480 50584 368532 50590
rect 368480 50526 368532 50532
rect 361580 46436 361632 46442
rect 361580 46378 361632 46384
rect 361592 16574 361620 46378
rect 365720 42288 365772 42294
rect 365720 42230 365772 42236
rect 362960 36780 363012 36786
rect 362960 36722 363012 36728
rect 362972 16574 363000 36722
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 361120 14748 361172 14754
rect 361120 14690 361172 14696
rect 357532 10600 357584 10606
rect 357532 10542 357584 10548
rect 357544 3602 357572 10542
rect 359924 7744 359976 7750
rect 359924 7686 359976 7692
rect 357532 3596 357584 3602
rect 357532 3538 357584 3544
rect 358728 3596 358780 3602
rect 358728 3538 358780 3544
rect 357452 3454 357572 3482
rect 357544 480 357572 3454
rect 358740 480 358768 3538
rect 359936 480 359964 7686
rect 361132 480 361160 14690
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364616 14680 364668 14686
rect 364616 14622 364668 14628
rect 364628 480 364656 14622
rect 365732 3482 365760 42230
rect 365812 36712 365864 36718
rect 365812 36654 365864 36660
rect 365824 3602 365852 36654
rect 368492 16574 368520 50526
rect 369860 45008 369912 45014
rect 369860 44950 369912 44956
rect 369872 16574 369900 44950
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 367744 14612 367796 14618
rect 367744 14554 367796 14560
rect 365812 3596 365864 3602
rect 365812 3538 365864 3544
rect 367008 3596 367060 3602
rect 367008 3538 367060 3544
rect 365732 3454 365852 3482
rect 365824 480 365852 3454
rect 367020 480 367048 3538
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 14554
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 66982
rect 372620 61464 372672 61470
rect 372620 61406 372672 61412
rect 372632 16574 372660 61406
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3602 374040 75346
rect 378140 72684 378192 72690
rect 378140 72626 378192 72632
rect 376760 46368 376812 46374
rect 376760 46310 376812 46316
rect 374092 38208 374144 38214
rect 374092 38150 374144 38156
rect 374000 3596 374052 3602
rect 374000 3538 374052 3544
rect 374104 480 374132 38150
rect 375380 29844 375432 29850
rect 375380 29786 375432 29792
rect 375392 16574 375420 29786
rect 376772 16574 376800 46310
rect 378152 16574 378180 72626
rect 382280 69896 382332 69902
rect 382280 69838 382332 69844
rect 380900 38140 380952 38146
rect 380900 38082 380952 38088
rect 379520 27124 379572 27130
rect 379520 27066 379572 27072
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 375288 3596 375340 3602
rect 375288 3538 375340 3544
rect 375300 480 375328 3538
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 27066
rect 380912 16574 380940 38082
rect 382292 16574 382320 69838
rect 398840 69828 398892 69834
rect 398840 69770 398892 69776
rect 385040 68536 385092 68542
rect 385040 68478 385092 68484
rect 383660 38072 383712 38078
rect 383660 38014 383712 38020
rect 383672 16574 383700 38014
rect 385052 16574 385080 68478
rect 391940 68468 391992 68474
rect 391940 68410 391992 68416
rect 389180 66972 389232 66978
rect 389180 66914 389232 66920
rect 387800 39636 387852 39642
rect 387800 39578 387852 39584
rect 380912 16546 381216 16574
rect 382292 16546 382412 16574
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 381188 480 381216 16546
rect 382384 480 382412 16546
rect 383568 6316 383620 6322
rect 383568 6258 383620 6264
rect 383580 480 383608 6258
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 387156 9240 387208 9246
rect 387156 9182 387208 9188
rect 387168 480 387196 9182
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 354 387840 39578
rect 389192 16574 389220 66914
rect 390560 39568 390612 39574
rect 390560 39510 390612 39516
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3602 390600 39510
rect 391952 16574 391980 68410
rect 396080 68400 396132 68406
rect 396080 68342 396132 68348
rect 391952 16546 392624 16574
rect 390652 14544 390704 14550
rect 390652 14486 390704 14492
rect 390560 3596 390612 3602
rect 390560 3538 390612 3544
rect 390664 480 390692 14486
rect 391848 3596 391900 3602
rect 391848 3538 391900 3544
rect 391860 480 391888 3538
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 395344 9172 395396 9178
rect 395344 9114 395396 9120
rect 394240 7676 394292 7682
rect 394240 7618 394292 7624
rect 394252 480 394280 7618
rect 395356 480 395384 9114
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 68342
rect 397460 19984 397512 19990
rect 397460 19926 397512 19932
rect 397472 16574 397500 19926
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3602 398880 69770
rect 402980 69760 403032 69766
rect 402980 69702 403032 69708
rect 398932 40928 398984 40934
rect 398932 40870 398984 40876
rect 398840 3596 398892 3602
rect 398840 3538 398892 3544
rect 398944 480 398972 40870
rect 400220 39500 400272 39506
rect 400220 39442 400272 39448
rect 400232 16574 400260 39442
rect 401600 39432 401652 39438
rect 401600 39374 401652 39380
rect 401612 16574 401640 39374
rect 402992 16574 403020 69702
rect 405740 46300 405792 46306
rect 405740 46242 405792 46248
rect 404360 21412 404412 21418
rect 404360 21354 404412 21360
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 400128 3596 400180 3602
rect 400128 3538 400180 3544
rect 400140 480 400168 3538
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 21354
rect 405752 16574 405780 46242
rect 407120 31136 407172 31142
rect 407120 31078 407172 31084
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 2650 407160 31078
rect 407212 16108 407264 16114
rect 407212 16050 407264 16056
rect 407120 2644 407172 2650
rect 407120 2586 407172 2592
rect 407224 480 407252 16050
rect 407776 3806 407804 77998
rect 411904 77988 411956 77994
rect 411904 77930 411956 77936
rect 411260 32496 411312 32502
rect 411260 32438 411312 32444
rect 410800 16040 410852 16046
rect 410800 15982 410852 15988
rect 409604 9104 409656 9110
rect 409604 9046 409656 9052
rect 407764 3800 407816 3806
rect 407764 3742 407816 3748
rect 408408 2644 408460 2650
rect 408408 2586 408460 2592
rect 408420 480 408448 2586
rect 409616 480 409644 9046
rect 410812 480 410840 15982
rect 411272 6914 411300 32438
rect 411916 16574 411944 77930
rect 414020 71256 414072 71262
rect 414020 71198 414072 71204
rect 412640 46232 412692 46238
rect 412640 46174 412692 46180
rect 411916 16546 412036 16574
rect 411272 6886 411944 6914
rect 411916 480 411944 6886
rect 412008 3738 412036 16546
rect 411996 3732 412048 3738
rect 411996 3674 412048 3680
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 46174
rect 414032 16574 414060 71198
rect 415400 42220 415452 42226
rect 415400 42162 415452 42168
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 2922 415440 42162
rect 418160 36644 418212 36650
rect 418160 36586 418212 36592
rect 415492 33856 415544 33862
rect 415492 33798 415544 33804
rect 415400 2916 415452 2922
rect 415400 2858 415452 2864
rect 415504 480 415532 33798
rect 418172 16574 418200 36586
rect 418172 16546 418568 16574
rect 417424 15972 417476 15978
rect 417424 15914 417476 15920
rect 416688 2916 416740 2922
rect 416688 2858 416740 2864
rect 416700 480 416728 2858
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 15914
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 418816 3602 418844 78134
rect 422944 78124 422996 78130
rect 422944 78066 422996 78072
rect 420920 71188 420972 71194
rect 420920 71130 420972 71136
rect 419540 42152 419592 42158
rect 419540 42094 419592 42100
rect 419552 16574 419580 42094
rect 419552 16546 420224 16574
rect 418804 3596 418856 3602
rect 418804 3538 418856 3544
rect 420196 480 420224 16546
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 71130
rect 422300 38004 422352 38010
rect 422300 37946 422352 37952
rect 422312 16574 422340 37946
rect 422312 16546 422616 16574
rect 422588 480 422616 16546
rect 422956 3670 422984 78066
rect 441620 76764 441672 76770
rect 441620 76706 441672 76712
rect 434720 75336 434772 75342
rect 434720 75278 434772 75284
rect 431960 74044 432012 74050
rect 431960 73986 432012 73992
rect 427820 72616 427872 72622
rect 427820 72558 427872 72564
rect 423680 71120 423732 71126
rect 423680 71062 423732 71068
rect 422944 3664 422996 3670
rect 422944 3606 422996 3612
rect 423692 3398 423720 71062
rect 425060 44940 425112 44946
rect 425060 44882 425112 44888
rect 425072 16574 425100 44882
rect 426440 43716 426492 43722
rect 426440 43658 426492 43664
rect 426452 16574 426480 43658
rect 427832 16574 427860 72558
rect 430580 43580 430632 43586
rect 430580 43522 430632 43528
rect 429200 24404 429252 24410
rect 429200 24346 429252 24352
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 423772 9036 423824 9042
rect 423772 8978 423824 8984
rect 423680 3392 423732 3398
rect 423680 3334 423732 3340
rect 423784 480 423812 8978
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 24346
rect 430592 16574 430620 43522
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 1170 432000 73986
rect 432052 43648 432104 43654
rect 432052 43590 432104 43596
rect 432064 3398 432092 43590
rect 433340 43512 433392 43518
rect 433340 43454 433392 43460
rect 433352 16574 433380 43454
rect 434732 16574 434760 75278
rect 438860 75268 438912 75274
rect 438860 75210 438912 75216
rect 436100 53304 436152 53310
rect 436100 53246 436152 53252
rect 436112 16574 436140 53246
rect 438872 16574 438900 75210
rect 440332 47864 440384 47870
rect 440332 47806 440384 47812
rect 440240 47796 440292 47802
rect 440240 47738 440292 47744
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 438872 16546 439176 16574
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 431972 1142 432092 1170
rect 432064 480 432092 1142
rect 433260 480 433288 3334
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 437940 5024 437992 5030
rect 437940 4966 437992 4972
rect 437952 480 437980 4966
rect 439148 480 439176 16546
rect 440252 3398 440280 47738
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 47806
rect 441632 16574 441660 76706
rect 445760 76696 445812 76702
rect 445760 76638 445812 76644
rect 444380 47728 444432 47734
rect 444380 47670 444432 47676
rect 443000 40860 443052 40866
rect 443000 40802 443052 40808
rect 443012 16574 443040 40802
rect 444392 16574 444420 47670
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 76638
rect 469220 76628 469272 76634
rect 469220 76570 469272 76576
rect 465080 57452 465132 57458
rect 465080 57394 465132 57400
rect 456800 56092 456852 56098
rect 456800 56034 456852 56040
rect 447140 54800 447192 54806
rect 447140 54742 447192 54748
rect 447152 16574 447180 54742
rect 451280 49156 451332 49162
rect 451280 49098 451332 49104
rect 448520 47660 448572 47666
rect 448520 47602 448572 47608
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 3210 448560 47602
rect 448612 32428 448664 32434
rect 448612 32370 448664 32376
rect 448624 3398 448652 32370
rect 449900 22908 449952 22914
rect 449900 22850 449952 22856
rect 449912 16574 449940 22850
rect 451292 16574 451320 49098
rect 455420 49088 455472 49094
rect 455420 49030 455472 49036
rect 455432 16574 455460 49030
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 455432 16546 455736 16574
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 454040 13320 454092 13326
rect 454040 13262 454092 13268
rect 453304 8968 453356 8974
rect 453304 8910 453356 8916
rect 453316 480 453344 8910
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 13262
rect 455708 480 455736 16546
rect 456812 3398 456840 56034
rect 462320 50516 462372 50522
rect 462320 50458 462372 50464
rect 458180 49020 458232 49026
rect 458180 48962 458232 48968
rect 458192 16574 458220 48962
rect 458192 16546 459232 16574
rect 456892 10532 456944 10538
rect 456892 10474 456944 10480
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 10474
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 459928 13252 459980 13258
rect 459928 13194 459980 13200
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 13194
rect 461584 3800 461636 3806
rect 461584 3742 461636 3748
rect 461596 480 461624 3742
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 50458
rect 463976 14476 464028 14482
rect 463976 14418 464028 14424
rect 463988 480 464016 14418
rect 465092 6914 465120 57394
rect 465172 50448 465224 50454
rect 465172 50390 465224 50396
rect 465184 16574 465212 50390
rect 469232 16574 469260 76570
rect 546500 75200 546552 75206
rect 546500 75142 546552 75148
rect 514760 73976 514812 73982
rect 514760 73918 514812 73924
rect 485780 61396 485832 61402
rect 485780 61338 485832 61344
rect 471980 58880 472032 58886
rect 471980 58822 472032 58828
rect 470600 31068 470652 31074
rect 470600 31010 470652 31016
rect 465184 16546 465856 16574
rect 469232 16546 469904 16574
rect 465092 6886 465212 6914
rect 465184 480 465212 6886
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467472 15904 467524 15910
rect 467472 15846 467524 15852
rect 467484 480 467512 15846
rect 468668 3732 468720 3738
rect 468668 3674 468720 3680
rect 468680 480 468708 3674
rect 469876 480 469904 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 31010
rect 471992 16574 472020 58822
rect 476120 51876 476172 51882
rect 476120 51818 476172 51824
rect 473360 50380 473412 50386
rect 473360 50322 473412 50328
rect 473372 16574 473400 50322
rect 476132 16574 476160 51818
rect 481640 44872 481692 44878
rect 481640 44814 481692 44820
rect 477500 33788 477552 33794
rect 477500 33730 477552 33736
rect 477512 16574 477540 33730
rect 480260 22840 480312 22846
rect 480260 22782 480312 22788
rect 480272 16574 480300 22782
rect 471992 16546 472296 16574
rect 473372 16546 473492 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 472268 480 472296 16546
rect 473464 480 473492 16546
rect 474096 13184 474148 13190
rect 474096 13126 474148 13132
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 13126
rect 475752 6248 475804 6254
rect 475752 6190 475804 6196
rect 475764 480 475792 6190
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 481652 3534 481680 44814
rect 483020 42084 483072 42090
rect 483020 42026 483072 42032
rect 483032 16574 483060 42026
rect 485792 16574 485820 61338
rect 509240 54732 509292 54738
rect 509240 54674 509292 54680
rect 498200 53236 498252 53242
rect 498200 53178 498252 53184
rect 491300 51808 491352 51814
rect 491300 51750 491352 51756
rect 487160 24336 487212 24342
rect 487160 24278 487212 24284
rect 483032 16546 484072 16574
rect 485792 16546 486464 16574
rect 481732 10464 481784 10470
rect 481732 10406 481784 10412
rect 481640 3528 481692 3534
rect 481640 3470 481692 3476
rect 481744 480 481772 10406
rect 482468 3528 482520 3534
rect 482468 3470 482520 3476
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3470
rect 484044 480 484072 16546
rect 484768 10396 484820 10402
rect 484768 10338 484820 10344
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 10338
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 24278
rect 489920 24268 489972 24274
rect 489920 24210 489972 24216
rect 488816 10328 488868 10334
rect 488816 10270 488868 10276
rect 488828 480 488856 10270
rect 489932 3534 489960 24210
rect 491312 16574 491340 51750
rect 495440 51740 495492 51746
rect 495440 51682 495492 51688
rect 494060 24200 494112 24206
rect 494060 24142 494112 24148
rect 492680 17468 492732 17474
rect 492680 17410 492732 17416
rect 492692 16574 492720 17410
rect 494072 16574 494100 24142
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 490012 11960 490064 11966
rect 490012 11902 490064 11908
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 11902
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 51682
rect 496820 17400 496872 17406
rect 496820 17342 496872 17348
rect 496832 16574 496860 17342
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 3534 498240 53178
rect 502340 53168 502392 53174
rect 502340 53110 502392 53116
rect 498292 25696 498344 25702
rect 498292 25638 498344 25644
rect 498200 3528 498252 3534
rect 498200 3470 498252 3476
rect 498304 3346 498332 25638
rect 500960 25628 501012 25634
rect 500960 25570 501012 25576
rect 499580 17332 499632 17338
rect 499580 17274 499632 17280
rect 499592 16574 499620 17274
rect 500972 16574 501000 25570
rect 502352 16574 502380 53110
rect 506480 53100 506532 53106
rect 506480 53042 506532 53048
rect 505100 43444 505152 43450
rect 505100 43386 505152 43392
rect 503720 17264 503772 17270
rect 503720 17206 503772 17212
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 499028 3528 499080 3534
rect 499028 3470 499080 3476
rect 498212 3318 498332 3346
rect 498212 480 498240 3318
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3470
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 17206
rect 505112 16574 505140 43386
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 480 506520 53042
rect 506572 36576 506624 36582
rect 506572 36518 506624 36524
rect 506584 16574 506612 36518
rect 507860 25560 507912 25566
rect 507860 25502 507912 25508
rect 507872 16574 507900 25502
rect 509252 16574 509280 54674
rect 513380 54664 513432 54670
rect 513380 54606 513432 54612
rect 510620 37936 510672 37942
rect 510620 37878 510672 37884
rect 510632 16574 510660 37878
rect 512000 27056 512052 27062
rect 512000 26998 512052 27004
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 26998
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 54606
rect 514772 3534 514800 73918
rect 527180 73908 527232 73914
rect 527180 73850 527232 73856
rect 517520 64184 517572 64190
rect 517520 64126 517572 64132
rect 514852 62824 514904 62830
rect 514852 62766 514904 62772
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 62766
rect 516140 54596 516192 54602
rect 516140 54538 516192 54544
rect 516152 16574 516180 54538
rect 517532 16574 517560 64126
rect 520280 56024 520332 56030
rect 520280 55966 520332 55972
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 5024 519596 5030
rect 519544 4966 519596 4972
rect 519556 480 519584 4966
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 55966
rect 523040 55956 523092 55962
rect 523040 55898 523092 55904
rect 521660 22772 521712 22778
rect 521660 22714 521712 22720
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 22714
rect 523052 3534 523080 55898
rect 523132 26988 523184 26994
rect 523132 26930 523184 26936
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523144 3346 523172 26930
rect 525800 26920 525852 26926
rect 525800 26862 525852 26868
rect 524420 24132 524472 24138
rect 524420 24074 524472 24080
rect 524432 16574 524460 24074
rect 525812 16574 525840 26862
rect 527192 16574 527220 73850
rect 540980 73840 541032 73846
rect 540980 73782 541032 73788
rect 529940 72548 529992 72554
rect 529940 72490 529992 72496
rect 528560 40792 528612 40798
rect 528560 40734 528612 40740
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 523868 3528 523920 3534
rect 523868 3470 523920 3476
rect 523052 3318 523172 3346
rect 523052 480 523080 3318
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523880 354 523908 3470
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 40734
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 72490
rect 539600 72480 539652 72486
rect 539600 72422 539652 72428
rect 534080 57384 534132 57390
rect 534080 57326 534132 57332
rect 531320 55888 531372 55894
rect 531320 55830 531372 55836
rect 531332 480 531360 55830
rect 531412 39364 531464 39370
rect 531412 39306 531464 39312
rect 531424 16574 531452 39306
rect 532700 28416 532752 28422
rect 532700 28358 532752 28364
rect 532712 16574 532740 28358
rect 534092 16574 534120 57326
rect 538220 57316 538272 57322
rect 538220 57258 538272 57264
rect 535460 47592 535512 47598
rect 535460 47534 535512 47540
rect 535472 16574 535500 47534
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537208 4888 537260 4894
rect 537208 4830 537260 4836
rect 537220 480 537248 4830
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 57258
rect 539612 3534 539640 72422
rect 539692 18828 539744 18834
rect 539692 18770 539744 18776
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 18770
rect 540992 16574 541020 73782
rect 542360 65544 542412 65550
rect 542360 65486 542412 65492
rect 542372 16574 542400 65486
rect 543740 60104 543792 60110
rect 543740 60046 543792 60052
rect 543752 16574 543780 60046
rect 545120 57248 545172 57254
rect 545120 57190 545172 57196
rect 545132 16574 545160 57190
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 75142
rect 556160 68332 556212 68338
rect 556160 68274 556212 68280
rect 553400 66904 553452 66910
rect 553400 66846 553452 66852
rect 550088 46912 550140 46918
rect 550086 46880 550088 46889
rect 550548 46912 550600 46918
rect 550140 46880 550142 46889
rect 550548 46854 550600 46860
rect 550086 46815 550142 46824
rect 550560 46238 550588 46854
rect 550548 46232 550600 46238
rect 550548 46174 550600 46180
rect 550640 28348 550692 28354
rect 550640 28290 550692 28296
rect 550652 16574 550680 28290
rect 553412 16574 553440 66846
rect 554780 28280 554832 28286
rect 554780 28222 554832 28228
rect 550652 16546 551048 16574
rect 553412 16546 553808 16574
rect 550272 13116 550324 13122
rect 550272 13058 550324 13064
rect 548616 11892 548668 11898
rect 548616 11834 548668 11840
rect 547880 4820 547932 4826
rect 547880 4762 547932 4768
rect 547892 480 547920 4762
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 11834
rect 550284 480 550312 13058
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552664 11824 552716 11830
rect 552664 11766 552716 11772
rect 552676 480 552704 11766
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 28222
rect 556172 3534 556200 68274
rect 559012 40724 559064 40730
rect 559012 40666 559064 40672
rect 557540 29776 557592 29782
rect 557540 29718 557592 29724
rect 557552 16574 557580 29718
rect 559024 16574 559052 40666
rect 560128 20670 560156 420022
rect 560220 419830 560248 420951
rect 560298 420472 560354 420481
rect 560298 420407 560354 420416
rect 560208 419824 560260 419830
rect 560208 419766 560260 419772
rect 560312 86902 560340 420407
rect 560392 420028 560444 420034
rect 560392 419970 560444 419976
rect 560404 167006 560432 419970
rect 560496 206990 560524 421087
rect 560588 245614 560616 421223
rect 560680 298790 560708 421806
rect 560760 421796 560812 421802
rect 560760 421738 560812 421744
rect 560772 353258 560800 421738
rect 560944 421320 560996 421326
rect 560944 421262 560996 421268
rect 560760 353252 560812 353258
rect 560760 353194 560812 353200
rect 560772 352578 560800 353194
rect 560760 352572 560812 352578
rect 560760 352514 560812 352520
rect 560668 298784 560720 298790
rect 560668 298726 560720 298732
rect 560576 245608 560628 245614
rect 560576 245550 560628 245556
rect 560588 244934 560616 245550
rect 560576 244928 560628 244934
rect 560576 244870 560628 244876
rect 560484 206984 560536 206990
rect 560484 206926 560536 206932
rect 560496 206310 560524 206926
rect 560484 206304 560536 206310
rect 560484 206246 560536 206252
rect 560392 167000 560444 167006
rect 560392 166942 560444 166948
rect 560300 86896 560352 86902
rect 560300 86838 560352 86844
rect 560956 20670 560984 421262
rect 561048 60722 561076 422758
rect 561680 422612 561732 422618
rect 561680 422554 561732 422560
rect 561128 421252 561180 421258
rect 561128 421194 561180 421200
rect 561140 73166 561168 421194
rect 561220 421116 561272 421122
rect 561220 421058 561272 421064
rect 561232 113150 561260 421058
rect 561692 419490 561720 422554
rect 580816 421932 580868 421938
rect 580816 421874 580868 421880
rect 580724 421728 580776 421734
rect 580724 421670 580776 421676
rect 580540 421660 580592 421666
rect 580540 421602 580592 421608
rect 563888 421524 563940 421530
rect 563888 421466 563940 421472
rect 563796 421456 563848 421462
rect 563796 421398 563848 421404
rect 562416 421388 562468 421394
rect 562416 421330 562468 421336
rect 562324 421048 562376 421054
rect 562324 420990 562376 420996
rect 561680 419484 561732 419490
rect 561680 419426 561732 419432
rect 561678 418568 561734 418577
rect 561678 418503 561734 418512
rect 561588 299464 561640 299470
rect 561588 299406 561640 299412
rect 561600 298790 561628 299406
rect 561588 298784 561640 298790
rect 561588 298726 561640 298732
rect 561312 201476 561364 201482
rect 561312 201418 561364 201424
rect 561324 200190 561352 201418
rect 561312 200184 561364 200190
rect 561312 200126 561364 200132
rect 561220 113144 561272 113150
rect 561220 113086 561272 113092
rect 561128 73160 561180 73166
rect 561128 73102 561180 73108
rect 561036 60716 561088 60722
rect 561036 60658 561088 60664
rect 560116 20664 560168 20670
rect 560116 20606 560168 20612
rect 560944 20664 560996 20670
rect 560944 20606 560996 20612
rect 560300 18760 560352 18766
rect 560300 18702 560352 18708
rect 560312 16574 560340 18702
rect 557552 16546 558592 16574
rect 559024 16546 559328 16574
rect 560312 16546 560432 16574
rect 556252 11756 556304 11762
rect 556252 11698 556304 11704
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556264 3346 556292 11698
rect 556988 3528 557040 3534
rect 556988 3470 557040 3476
rect 556172 3318 556292 3346
rect 556172 480 556200 3318
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557000 354 557028 3470
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 561324 6866 561352 200126
rect 561692 7614 561720 418503
rect 561770 416120 561826 416129
rect 561770 416055 561826 416064
rect 561680 7608 561732 7614
rect 561680 7550 561732 7556
rect 561312 6860 561364 6866
rect 561312 6802 561364 6808
rect 561784 6186 561812 416055
rect 562336 193186 562364 420990
rect 562428 273222 562456 421330
rect 562508 420096 562560 420102
rect 562508 420038 562560 420044
rect 562520 405686 562548 420038
rect 563704 419620 563756 419626
rect 563704 419562 563756 419568
rect 562508 405680 562560 405686
rect 562508 405622 562560 405628
rect 562416 273216 562468 273222
rect 562416 273158 562468 273164
rect 563716 259418 563744 419562
rect 563808 325650 563836 421398
rect 563900 379506 563928 421466
rect 580264 421184 580316 421190
rect 580264 421126 580316 421132
rect 569224 420980 569276 420986
rect 569224 420922 569276 420928
rect 566464 419552 566516 419558
rect 566464 419494 566516 419500
rect 563888 379500 563940 379506
rect 563888 379442 563940 379448
rect 564438 371920 564494 371929
rect 564438 371855 564494 371864
rect 563796 325644 563848 325650
rect 563796 325586 563848 325592
rect 563704 259412 563756 259418
rect 563704 259354 563756 259360
rect 564452 201482 564480 371855
rect 566476 313274 566504 419494
rect 566464 313268 566516 313274
rect 566464 313210 566516 313216
rect 564440 201476 564492 201482
rect 564440 201418 564492 201424
rect 562324 193180 562376 193186
rect 562324 193122 562376 193128
rect 569236 179382 569264 420922
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 579620 353252 579672 353258
rect 579620 353194 579672 353200
rect 579632 351937 579660 353194
rect 579618 351928 579674 351937
rect 579618 351863 579674 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 579620 193180 579672 193186
rect 579620 193122 579672 193128
rect 579632 192545 579660 193122
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 569224 179376 569276 179382
rect 569224 179318 569276 179324
rect 579620 179376 579672 179382
rect 579620 179318 579672 179324
rect 579632 179217 579660 179318
rect 579618 179208 579674 179217
rect 579618 179143 579674 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579620 113144 579672 113150
rect 579620 113086 579672 113092
rect 579632 112849 579660 113086
rect 579618 112840 579674 112849
rect 579618 112775 579674 112784
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 574100 76560 574152 76566
rect 574100 76502 574152 76508
rect 571340 71052 571392 71058
rect 571340 70994 571392 71000
rect 564532 69692 564584 69698
rect 564532 69634 564584 69640
rect 563060 58812 563112 58818
rect 563060 58754 563112 58760
rect 561864 29708 561916 29714
rect 561864 29650 561916 29656
rect 561876 16574 561904 29650
rect 561876 16546 562088 16574
rect 561772 6180 561824 6186
rect 561772 6122 561824 6128
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 58754
rect 564544 6914 564572 69634
rect 565820 58744 565872 58750
rect 565820 58686 565872 58692
rect 564624 35352 564676 35358
rect 564624 35294 564676 35300
rect 564636 16574 564664 35294
rect 565832 16574 565860 58686
rect 569960 58676 570012 58682
rect 569960 58618 570012 58624
rect 568580 29640 568632 29646
rect 568580 29582 568632 29588
rect 567200 18692 567252 18698
rect 567200 18634 567252 18640
rect 567212 16574 567240 18634
rect 568592 16574 568620 29582
rect 569972 16574 570000 58618
rect 564636 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 564452 6886 564572 6914
rect 564452 480 564480 6886
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 70994
rect 572720 54528 572772 54534
rect 572720 54470 572772 54476
rect 572732 3534 572760 54470
rect 572812 35284 572864 35290
rect 572812 35226 572864 35232
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 572824 3346 572852 35226
rect 574112 16574 574140 76502
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 576860 60036 576912 60042
rect 576860 59978 576912 59984
rect 575480 35216 575532 35222
rect 575480 35158 575532 35164
rect 575492 16574 575520 35158
rect 576872 16574 576900 59978
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580184 46238 580212 46271
rect 580172 46232 580224 46238
rect 580172 46174 580224 46180
rect 580276 33153 580304 421126
rect 580356 420436 580408 420442
rect 580356 420378 580408 420384
rect 580368 99521 580396 420378
rect 580448 420368 580500 420374
rect 580448 420310 580500 420316
rect 580460 139369 580488 420310
rect 580552 152697 580580 421602
rect 580632 420300 580684 420306
rect 580632 420242 580684 420248
rect 580644 219065 580672 420242
rect 580736 232393 580764 421670
rect 580828 365129 580856 421874
rect 580814 365120 580870 365129
rect 580814 365055 580870 365064
rect 580722 232384 580778 232393
rect 580722 232319 580778 232328
rect 580630 219056 580686 219065
rect 580630 218991 580686 219000
rect 580538 152688 580594 152697
rect 580538 152623 580594 152632
rect 580446 139360 580502 139369
rect 580446 139295 580502 139304
rect 580354 99512 580410 99521
rect 580354 99447 580410 99456
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 578240 18624 578292 18630
rect 578240 18566 578292 18572
rect 578252 16574 578280 18566
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 573548 3528 573600 3534
rect 573548 3470 573600 3476
rect 572732 3318 572852 3346
rect 572732 480 572760 3318
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573560 354 573588 3470
rect 575124 480 575152 16546
rect 573886 354 573998 480
rect 573560 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 583392 3664 583444 3670
rect 583392 3606 583444 3612
rect 581000 3596 581052 3602
rect 581000 3538 581052 3544
rect 581012 480 581040 3538
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 583404 480 583432 3606
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632032 3478 632088
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3054 501744 3110 501800
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 475632 3570 475688
rect 3606 462576 3662 462632
rect 3698 449520 3754 449576
rect 4066 423544 4122 423600
rect 4802 423136 4858 423192
rect 3514 422456 3570 422512
rect 3422 421640 3478 421696
rect 3330 410488 3386 410544
rect 3330 371320 3386 371376
rect 3054 358400 3110 358456
rect 2962 345344 3018 345400
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3238 293120 3294 293176
rect 3330 267144 3386 267200
rect 2962 254088 3018 254144
rect 3330 214920 3386 214976
rect 2778 162832 2834 162888
rect 2778 149776 2834 149832
rect 2778 97552 2834 97608
rect 2962 84632 3018 84688
rect 3606 421776 3662 421832
rect 3514 188808 3570 188864
rect 3514 136720 3570 136776
rect 3790 421504 3846 421560
rect 3882 397432 3938 397488
rect 3790 241032 3846 241088
rect 3698 201864 3754 201920
rect 3698 71576 3754 71632
rect 3606 58520 3662 58576
rect 3422 45464 3478 45520
rect 3882 110608 3938 110664
rect 4986 422592 5042 422648
rect 79322 422728 79378 422784
rect 226982 419872 227038 419928
rect 223486 371220 223488 371240
rect 223488 371220 223540 371240
rect 223540 371220 223542 371240
rect 223486 371184 223542 371220
rect 444930 420280 444986 420336
rect 444746 420144 444802 420200
rect 445390 422864 445446 422920
rect 445574 420008 445630 420064
rect 3790 32408 3846 32464
rect 3422 19352 3478 19408
rect 142158 77424 142214 77480
rect 142526 77424 142582 77480
rect 169758 79872 169814 79928
rect 170264 79872 170320 79928
rect 521198 420416 521254 420472
rect 522394 420416 522450 420472
rect 523498 420960 523554 421016
rect 525614 421096 525670 421152
rect 527086 422320 527142 422376
rect 526626 421232 526682 421288
rect 535274 421776 535330 421832
rect 544014 422864 544070 422920
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580262 670656 580318 670712
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580354 564304 580410 564360
rect 580446 537784 580502 537840
rect 580538 511264 580594 511320
rect 551374 423000 551430 423056
rect 550638 421640 550694 421696
rect 552110 420144 552166 420200
rect 552754 420280 552810 420336
rect 552570 419872 552626 419928
rect 556158 422728 556214 422784
rect 553858 421504 553914 421560
rect 554870 422456 554926 422512
rect 555238 422320 555294 422376
rect 556342 422592 556398 422648
rect 557538 423136 557594 423192
rect 557814 420008 557870 420064
rect 560574 421232 560630 421288
rect 560482 421096 560538 421152
rect 560206 420960 560262 421016
rect 559194 419872 559250 419928
rect 517518 419600 517574 419656
rect 447598 365200 447654 365256
rect 447690 355408 447746 355464
rect 447874 367104 447930 367160
rect 447874 366424 447930 366480
rect 447782 345752 447838 345808
rect 447782 302912 447838 302968
rect 447966 326168 448022 326224
rect 448150 324264 448206 324320
rect 448058 322360 448114 322416
rect 448242 320456 448298 320512
rect 448334 318416 448390 318472
rect 448978 363160 449034 363216
rect 449070 361256 449126 361312
rect 449162 343712 449218 343768
rect 449346 341808 449402 341864
rect 449254 339904 449310 339960
rect 449530 337864 449586 337920
rect 449622 335960 449678 336016
rect 449438 334056 449494 334112
rect 449714 332016 449770 332072
rect 450726 369552 450782 369608
rect 450358 359896 450414 359952
rect 450266 357584 450322 357640
rect 450174 354048 450230 354104
rect 450082 351872 450138 351928
rect 449990 350104 450046 350160
rect 449898 347792 449954 347848
rect 449806 330112 449862 330168
rect 448426 316512 448482 316568
rect 447874 301008 447930 301064
rect 514022 385736 514078 385792
rect 514022 385056 514078 385112
rect 509974 384648 510030 384704
rect 510158 383968 510214 384024
rect 509974 383696 510030 383752
rect 510158 383696 510214 383752
rect 518162 419056 518218 419112
rect 517610 417832 517666 417888
rect 517518 416744 517574 416800
rect 517518 415520 517574 415576
rect 517518 414296 517574 414352
rect 517518 413208 517574 413264
rect 517518 411984 517574 412040
rect 517794 411440 517850 411496
rect 517518 410760 517574 410816
rect 517518 409672 517574 409728
rect 517610 408448 517666 408504
rect 517518 407244 517574 407280
rect 517518 407224 517520 407244
rect 517520 407224 517572 407244
rect 517572 407224 517574 407244
rect 517518 406136 517574 406192
rect 517518 404912 517574 404968
rect 517886 407904 517942 407960
rect 517702 403688 517758 403744
rect 517702 402600 517758 402656
rect 517794 401376 517850 401432
rect 517702 400308 517758 400344
rect 517702 400288 517704 400308
rect 517704 400288 517756 400308
rect 517756 400288 517758 400308
rect 517702 399064 517758 399120
rect 517702 397840 517758 397896
rect 517702 396752 517758 396808
rect 517886 396072 517942 396128
rect 517794 395528 517850 395584
rect 517702 394984 517758 395040
rect 517702 393760 517758 393816
rect 517702 391992 517758 392048
rect 517702 390768 517758 390824
rect 517702 389680 517758 389736
rect 517702 387932 517758 387968
rect 517702 387912 517704 387932
rect 517704 387912 517756 387932
rect 517756 387912 517758 387932
rect 517702 386688 517758 386744
rect 517886 393216 517942 393272
rect 517978 392536 518034 392592
rect 517886 391448 517942 391504
rect 517886 390224 517942 390280
rect 517978 389000 518034 389056
rect 517886 388456 517942 388512
rect 517886 387232 517942 387288
rect 518070 380840 518126 380896
rect 517794 378936 517850 378992
rect 518070 372000 518126 372056
rect 519910 419328 519966 419384
rect 518806 417288 518862 417344
rect 518714 416064 518770 416120
rect 518622 414976 518678 415032
rect 518530 413752 518586 413808
rect 518346 412528 518402 412584
rect 518254 410216 518310 410272
rect 518530 370912 518586 370968
rect 518346 370640 518402 370696
rect 518898 408992 518954 409048
rect 518990 406680 519046 406736
rect 519266 405456 519322 405512
rect 519082 404368 519138 404424
rect 519174 403144 519230 403200
rect 519358 401920 519414 401976
rect 519450 400832 519506 400888
rect 519542 399608 519598 399664
rect 519726 398520 519782 398576
rect 519542 379072 519598 379128
rect 519726 378800 519782 378856
rect 549350 315696 549406 315752
rect 549350 307128 549406 307184
rect 451462 299512 451518 299568
rect 454498 297880 454554 297936
rect 457626 297744 457682 297800
rect 488906 297880 488962 297936
rect 492034 297744 492090 297800
rect 495162 297608 495218 297664
rect 485778 297200 485834 297256
rect 548614 298016 548670 298072
rect 532698 297472 532754 297528
rect 529570 297336 529626 297392
rect 549902 363840 549958 363896
rect 550086 367784 550142 367840
rect 550086 350376 550142 350432
rect 551466 359080 551522 359136
rect 551374 354728 551430 354784
rect 551282 345888 551338 345944
rect 553398 370504 553454 370560
rect 552478 341536 552534 341592
rect 552386 337184 552442 337240
rect 552294 332832 552350 332888
rect 552202 328480 552258 328536
rect 552110 323992 552166 324048
rect 552018 319640 552074 319696
rect 551190 310936 551246 310992
rect 551098 302232 551154 302288
rect 553766 298016 553822 298072
rect 550086 46860 550088 46880
rect 550088 46860 550140 46880
rect 550140 46860 550142 46880
rect 550086 46824 550142 46860
rect 560298 420416 560354 420472
rect 561678 418512 561734 418568
rect 561770 416064 561826 416120
rect 564438 371864 564494 371920
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579618 351872 579674 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579802 205672 579858 205728
rect 579618 192480 579674 192536
rect 579618 179152 579674 179208
rect 580170 165824 580226 165880
rect 580170 125976 580226 126032
rect 579618 112784 579674 112840
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580814 365064 580870 365120
rect 580722 232328 580778 232384
rect 580630 219000 580686 219056
rect 580538 152632 580594 152688
rect 580446 139304 580502 139360
rect 580354 99456 580410 99512
rect 580262 33088 580318 33144
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 580349 564362 580415 564365
rect 583520 564362 584960 564452
rect 580349 564360 584960 564362
rect 580349 564304 580354 564360
rect 580410 564304 584960 564360
rect 580349 564302 584960 564304
rect 580349 564299 580415 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580441 537842 580507 537845
rect 583520 537842 584960 537932
rect 580441 537840 584960 537842
rect 580441 537784 580446 537840
rect 580502 537784 584960 537840
rect 580441 537782 584960 537784
rect 580441 537779 580507 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580533 511322 580599 511325
rect 583520 511322 584960 511412
rect 580533 511320 584960 511322
rect 580533 511264 580538 511320
rect 580594 511264 584960 511320
rect 580533 511262 584960 511264
rect 580533 511259 580599 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3509 475690 3575 475693
rect -960 475688 3575 475690
rect -960 475632 3514 475688
rect 3570 475632 3575 475688
rect -960 475630 3575 475632
rect -960 475540 480 475630
rect 3509 475627 3575 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3693 449578 3759 449581
rect -960 449576 3759 449578
rect -960 449520 3698 449576
rect 3754 449520 3759 449576
rect -960 449518 3759 449520
rect -960 449428 480 449518
rect 3693 449515 3759 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 4061 423602 4127 423605
rect -960 423600 4127 423602
rect -960 423544 4066 423600
rect 4122 423544 4127 423600
rect -960 423542 4127 423544
rect -960 423452 480 423542
rect 4061 423539 4127 423542
rect 4797 423194 4863 423197
rect 557533 423194 557599 423197
rect 4797 423192 557599 423194
rect 4797 423136 4802 423192
rect 4858 423136 557538 423192
rect 557594 423136 557599 423192
rect 4797 423134 557599 423136
rect 4797 423131 4863 423134
rect 557533 423131 557599 423134
rect 518014 422996 518020 423060
rect 518084 423058 518090 423060
rect 551369 423058 551435 423061
rect 518084 423056 551435 423058
rect 518084 423000 551374 423056
rect 551430 423000 551435 423056
rect 518084 422998 551435 423000
rect 518084 422996 518090 422998
rect 551369 422995 551435 422998
rect 445385 422922 445451 422925
rect 544009 422922 544075 422925
rect 445385 422920 544075 422922
rect 445385 422864 445390 422920
rect 445446 422864 544014 422920
rect 544070 422864 544075 422920
rect 445385 422862 544075 422864
rect 445385 422859 445451 422862
rect 544009 422859 544075 422862
rect 79317 422786 79383 422789
rect 556153 422786 556219 422789
rect 79317 422784 556219 422786
rect 79317 422728 79322 422784
rect 79378 422728 556158 422784
rect 556214 422728 556219 422784
rect 79317 422726 556219 422728
rect 79317 422723 79383 422726
rect 556153 422723 556219 422726
rect 4981 422650 5047 422653
rect 556337 422650 556403 422653
rect 4981 422648 556403 422650
rect 4981 422592 4986 422648
rect 5042 422592 556342 422648
rect 556398 422592 556403 422648
rect 4981 422590 556403 422592
rect 4981 422587 5047 422590
rect 556337 422587 556403 422590
rect 3509 422514 3575 422517
rect 554865 422514 554931 422517
rect 3509 422512 554931 422514
rect 3509 422456 3514 422512
rect 3570 422456 554870 422512
rect 554926 422456 554931 422512
rect 3509 422454 554931 422456
rect 3509 422451 3575 422454
rect 554865 422451 554931 422454
rect 527081 422378 527147 422381
rect 555233 422378 555299 422381
rect 527081 422376 555299 422378
rect 527081 422320 527086 422376
rect 527142 422320 555238 422376
rect 555294 422320 555299 422376
rect 527081 422318 555299 422320
rect 527081 422315 527147 422318
rect 555233 422315 555299 422318
rect 3601 421834 3667 421837
rect 535269 421834 535335 421837
rect 3601 421832 535335 421834
rect 3601 421776 3606 421832
rect 3662 421776 535274 421832
rect 535330 421776 535335 421832
rect 3601 421774 535335 421776
rect 3601 421771 3667 421774
rect 535269 421771 535335 421774
rect 3417 421698 3483 421701
rect 550633 421698 550699 421701
rect 3417 421696 550699 421698
rect 3417 421640 3422 421696
rect 3478 421640 550638 421696
rect 550694 421640 550699 421696
rect 3417 421638 550699 421640
rect 3417 421635 3483 421638
rect 550633 421635 550699 421638
rect 3785 421562 3851 421565
rect 553853 421562 553919 421565
rect 3785 421560 553919 421562
rect 3785 421504 3790 421560
rect 3846 421504 553858 421560
rect 553914 421504 553919 421560
rect 3785 421502 553919 421504
rect 3785 421499 3851 421502
rect 553853 421499 553919 421502
rect 526621 421290 526687 421293
rect 560569 421290 560635 421293
rect 526621 421288 560635 421290
rect 526621 421232 526626 421288
rect 526682 421232 560574 421288
rect 560630 421232 560635 421288
rect 526621 421230 560635 421232
rect 526621 421227 526687 421230
rect 560569 421227 560635 421230
rect 525609 421154 525675 421157
rect 560477 421154 560543 421157
rect 525609 421152 560543 421154
rect 525609 421096 525614 421152
rect 525670 421096 560482 421152
rect 560538 421096 560543 421152
rect 525609 421094 560543 421096
rect 525609 421091 525675 421094
rect 560477 421091 560543 421094
rect 523493 421018 523559 421021
rect 560201 421018 560267 421021
rect 523493 421016 560267 421018
rect 523493 420960 523498 421016
rect 523554 420960 560206 421016
rect 560262 420960 560267 421016
rect 523493 420958 560267 420960
rect 523493 420955 523559 420958
rect 560201 420955 560267 420958
rect 518750 420412 518756 420476
rect 518820 420474 518826 420476
rect 521193 420474 521259 420477
rect 518820 420472 521259 420474
rect 518820 420416 521198 420472
rect 521254 420416 521259 420472
rect 518820 420414 521259 420416
rect 518820 420412 518826 420414
rect 521193 420411 521259 420414
rect 522389 420474 522455 420477
rect 560293 420474 560359 420477
rect 522389 420472 560359 420474
rect 522389 420416 522394 420472
rect 522450 420416 560298 420472
rect 560354 420416 560359 420472
rect 522389 420414 560359 420416
rect 522389 420411 522455 420414
rect 560293 420411 560359 420414
rect 444925 420338 444991 420341
rect 552749 420338 552815 420341
rect 444925 420336 552815 420338
rect 444925 420280 444930 420336
rect 444986 420280 552754 420336
rect 552810 420280 552815 420336
rect 444925 420278 552815 420280
rect 444925 420275 444991 420278
rect 552749 420275 552815 420278
rect 444741 420202 444807 420205
rect 552105 420202 552171 420205
rect 444741 420200 552171 420202
rect 444741 420144 444746 420200
rect 444802 420144 552110 420200
rect 552166 420144 552171 420200
rect 444741 420142 552171 420144
rect 444741 420139 444807 420142
rect 552105 420139 552171 420142
rect 445569 420066 445635 420069
rect 557809 420066 557875 420069
rect 445569 420064 557875 420066
rect 445569 420008 445574 420064
rect 445630 420008 557814 420064
rect 557870 420008 557875 420064
rect 445569 420006 557875 420008
rect 445569 420003 445635 420006
rect 557809 420003 557875 420006
rect 226977 419930 227043 419933
rect 552565 419930 552631 419933
rect 226977 419928 552631 419930
rect 226977 419872 226982 419928
rect 227038 419872 552570 419928
rect 552626 419872 552631 419928
rect 226977 419870 552631 419872
rect 226977 419867 227043 419870
rect 552565 419867 552631 419870
rect 558862 419868 558868 419932
rect 558932 419930 558938 419932
rect 559189 419930 559255 419933
rect 558932 419928 559255 419930
rect 558932 419872 559194 419928
rect 559250 419872 559255 419928
rect 558932 419870 559255 419872
rect 558932 419868 558938 419870
rect 559189 419867 559255 419870
rect 517513 419658 517579 419661
rect 517513 419656 520076 419658
rect 517513 419600 517518 419656
rect 517574 419600 520076 419656
rect 517513 419598 520076 419600
rect 517513 419595 517579 419598
rect 519905 419388 519971 419389
rect 519854 419386 519860 419388
rect 519814 419326 519860 419386
rect 519924 419384 519971 419388
rect 519966 419328 519971 419384
rect 519854 419324 519860 419326
rect 519924 419324 519971 419328
rect 519905 419323 519971 419324
rect 518157 419114 518223 419117
rect 518157 419112 520076 419114
rect 518157 419056 518162 419112
rect 518218 419056 520076 419112
rect 518157 419054 520076 419056
rect 518157 419051 518223 419054
rect 518566 418508 518572 418572
rect 518636 418570 518642 418572
rect 559790 418570 559850 418812
rect 561673 418570 561739 418573
rect 518636 418510 520076 418570
rect 559790 418568 561739 418570
rect 559790 418512 561678 418568
rect 561734 418512 561739 418568
rect 559790 418510 561739 418512
rect 518636 418508 518642 418510
rect 561673 418507 561739 418510
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 517605 417890 517671 417893
rect 517605 417888 520076 417890
rect 517605 417832 517610 417888
rect 517666 417832 520076 417888
rect 517605 417830 520076 417832
rect 517605 417827 517671 417830
rect 518801 417346 518867 417349
rect 518801 417344 520076 417346
rect 518801 417288 518806 417344
rect 518862 417288 520076 417344
rect 518801 417286 520076 417288
rect 518801 417283 518867 417286
rect 517513 416802 517579 416805
rect 517513 416800 520076 416802
rect 517513 416744 517518 416800
rect 517574 416744 520076 416800
rect 517513 416742 520076 416744
rect 517513 416739 517579 416742
rect 518709 416122 518775 416125
rect 559790 416122 559850 416636
rect 561765 416122 561831 416125
rect 518709 416120 520076 416122
rect 518709 416064 518714 416120
rect 518770 416064 520076 416120
rect 518709 416062 520076 416064
rect 559790 416120 561831 416122
rect 559790 416064 561770 416120
rect 561826 416064 561831 416120
rect 559790 416062 561831 416064
rect 518709 416059 518775 416062
rect 561765 416059 561831 416062
rect 517513 415578 517579 415581
rect 517513 415576 520076 415578
rect 517513 415520 517518 415576
rect 517574 415520 520076 415576
rect 517513 415518 520076 415520
rect 517513 415515 517579 415518
rect 518617 415034 518683 415037
rect 518617 415032 520076 415034
rect 518617 414976 518622 415032
rect 518678 414976 520076 415032
rect 518617 414974 520076 414976
rect 518617 414971 518683 414974
rect 517513 414354 517579 414357
rect 517513 414352 520076 414354
rect 517513 414296 517518 414352
rect 517574 414296 520076 414352
rect 517513 414294 520076 414296
rect 517513 414291 517579 414294
rect 518525 413810 518591 413813
rect 518525 413808 520076 413810
rect 518525 413752 518530 413808
rect 518586 413752 520076 413808
rect 518525 413750 520076 413752
rect 518525 413747 518591 413750
rect 517513 413266 517579 413269
rect 517513 413264 520076 413266
rect 517513 413208 517518 413264
rect 517574 413208 520076 413264
rect 517513 413206 520076 413208
rect 517513 413203 517579 413206
rect 518341 412586 518407 412589
rect 518341 412584 520076 412586
rect 518341 412528 518346 412584
rect 518402 412528 520076 412584
rect 518341 412526 520076 412528
rect 518341 412523 518407 412526
rect 517513 412042 517579 412045
rect 517513 412040 520076 412042
rect 517513 411984 517518 412040
rect 517574 411984 520076 412040
rect 517513 411982 520076 411984
rect 517513 411979 517579 411982
rect 517789 411498 517855 411501
rect 517789 411496 520076 411498
rect 517789 411440 517794 411496
rect 517850 411440 520076 411496
rect 517789 411438 520076 411440
rect 517789 411435 517855 411438
rect 517513 410818 517579 410821
rect 517513 410816 520076 410818
rect 517513 410760 517518 410816
rect 517574 410760 520076 410816
rect 517513 410758 520076 410760
rect 517513 410755 517579 410758
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 518249 410274 518315 410277
rect 518249 410272 520076 410274
rect 518249 410216 518254 410272
rect 518310 410216 520076 410272
rect 518249 410214 520076 410216
rect 518249 410211 518315 410214
rect 517513 409730 517579 409733
rect 517513 409728 520076 409730
rect 517513 409672 517518 409728
rect 517574 409672 520076 409728
rect 517513 409670 520076 409672
rect 517513 409667 517579 409670
rect 518893 409050 518959 409053
rect 518893 409048 520076 409050
rect 518893 408992 518898 409048
rect 518954 408992 520076 409048
rect 518893 408990 520076 408992
rect 518893 408987 518959 408990
rect 517605 408506 517671 408509
rect 517605 408504 520076 408506
rect 517605 408448 517610 408504
rect 517666 408448 520076 408504
rect 517605 408446 520076 408448
rect 517605 408443 517671 408446
rect 517881 407962 517947 407965
rect 517881 407960 520076 407962
rect 517881 407904 517886 407960
rect 517942 407904 520076 407960
rect 517881 407902 520076 407904
rect 517881 407899 517947 407902
rect 517513 407282 517579 407285
rect 517513 407280 520076 407282
rect 517513 407224 517518 407280
rect 517574 407224 520076 407280
rect 517513 407222 520076 407224
rect 517513 407219 517579 407222
rect 518985 406738 519051 406741
rect 518985 406736 520076 406738
rect 518985 406680 518990 406736
rect 519046 406680 520076 406736
rect 518985 406678 520076 406680
rect 518985 406675 519051 406678
rect 517513 406194 517579 406197
rect 517513 406192 520076 406194
rect 517513 406136 517518 406192
rect 517574 406136 520076 406192
rect 517513 406134 520076 406136
rect 517513 406131 517579 406134
rect 519261 405514 519327 405517
rect 519261 405512 520076 405514
rect 519261 405456 519266 405512
rect 519322 405456 520076 405512
rect 519261 405454 520076 405456
rect 519261 405451 519327 405454
rect 517513 404970 517579 404973
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 517513 404968 520076 404970
rect 517513 404912 517518 404968
rect 517574 404912 520076 404968
rect 517513 404910 520076 404912
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 517513 404907 517579 404910
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 519077 404426 519143 404429
rect 519077 404424 520076 404426
rect 519077 404368 519082 404424
rect 519138 404368 520076 404424
rect 519077 404366 520076 404368
rect 519077 404363 519143 404366
rect 517697 403746 517763 403749
rect 517697 403744 520076 403746
rect 517697 403688 517702 403744
rect 517758 403688 520076 403744
rect 517697 403686 520076 403688
rect 517697 403683 517763 403686
rect 519169 403202 519235 403205
rect 519169 403200 520076 403202
rect 519169 403144 519174 403200
rect 519230 403144 520076 403200
rect 519169 403142 520076 403144
rect 519169 403139 519235 403142
rect 517697 402658 517763 402661
rect 517697 402656 520076 402658
rect 517697 402600 517702 402656
rect 517758 402600 520076 402656
rect 517697 402598 520076 402600
rect 517697 402595 517763 402598
rect 519353 401978 519419 401981
rect 519353 401976 520076 401978
rect 519353 401920 519358 401976
rect 519414 401920 520076 401976
rect 519353 401918 520076 401920
rect 519353 401915 519419 401918
rect 517789 401434 517855 401437
rect 517789 401432 520076 401434
rect 517789 401376 517794 401432
rect 517850 401376 520076 401432
rect 517789 401374 520076 401376
rect 517789 401371 517855 401374
rect 519445 400890 519511 400893
rect 519445 400888 520076 400890
rect 519445 400832 519450 400888
rect 519506 400832 520076 400888
rect 519445 400830 520076 400832
rect 519445 400827 519511 400830
rect 517697 400346 517763 400349
rect 517697 400344 520076 400346
rect 517697 400288 517702 400344
rect 517758 400288 520076 400344
rect 517697 400286 520076 400288
rect 517697 400283 517763 400286
rect 519537 399666 519603 399669
rect 519537 399664 520076 399666
rect 519537 399608 519542 399664
rect 519598 399608 520076 399664
rect 519537 399606 520076 399608
rect 519537 399603 519603 399606
rect 517697 399122 517763 399125
rect 517697 399120 520076 399122
rect 517697 399064 517702 399120
rect 517758 399064 520076 399120
rect 517697 399062 520076 399064
rect 517697 399059 517763 399062
rect 519721 398578 519787 398581
rect 519721 398576 520076 398578
rect 519721 398520 519726 398576
rect 519782 398520 520076 398576
rect 519721 398518 520076 398520
rect 519721 398515 519787 398518
rect 517697 397898 517763 397901
rect 517697 397896 520076 397898
rect 517697 397840 517702 397896
rect 517758 397840 520076 397896
rect 517697 397838 520076 397840
rect 517697 397835 517763 397838
rect -960 397490 480 397580
rect 3877 397490 3943 397493
rect -960 397488 3943 397490
rect -960 397432 3882 397488
rect 3938 397432 3943 397488
rect -960 397430 3943 397432
rect -960 397340 480 397430
rect 3877 397427 3943 397430
rect 518934 397292 518940 397356
rect 519004 397354 519010 397356
rect 519004 397294 520076 397354
rect 519004 397292 519010 397294
rect 517697 396810 517763 396813
rect 517697 396808 520076 396810
rect 517697 396752 517702 396808
rect 517758 396752 520076 396808
rect 517697 396750 520076 396752
rect 517697 396747 517763 396750
rect 517881 396130 517947 396133
rect 517881 396128 520076 396130
rect 517881 396072 517886 396128
rect 517942 396072 520076 396128
rect 517881 396070 520076 396072
rect 517881 396067 517947 396070
rect 517789 395586 517855 395589
rect 517789 395584 520076 395586
rect 517789 395528 517794 395584
rect 517850 395528 520076 395584
rect 517789 395526 520076 395528
rect 517789 395523 517855 395526
rect 517697 395042 517763 395045
rect 517697 395040 520076 395042
rect 517697 394984 517702 395040
rect 517758 394984 520076 395040
rect 517697 394982 520076 394984
rect 517697 394979 517763 394982
rect 520046 394090 520106 394332
rect 509190 394030 520106 394090
rect 449382 393484 449388 393548
rect 449452 393546 449458 393548
rect 509190 393546 509250 394030
rect 517697 393818 517763 393821
rect 517697 393816 520076 393818
rect 517697 393760 517702 393816
rect 517758 393760 520076 393816
rect 517697 393758 520076 393760
rect 517697 393755 517763 393758
rect 449452 393486 509250 393546
rect 449452 393484 449458 393486
rect 517881 393274 517947 393277
rect 517881 393272 520076 393274
rect 517881 393216 517886 393272
rect 517942 393216 520076 393272
rect 517881 393214 520076 393216
rect 517881 393211 517947 393214
rect 517973 392594 518039 392597
rect 517973 392592 520076 392594
rect 517973 392536 517978 392592
rect 518034 392536 520076 392592
rect 517973 392534 520076 392536
rect 517973 392531 518039 392534
rect 517697 392050 517763 392053
rect 517697 392048 520076 392050
rect 517697 391992 517702 392048
rect 517758 391992 520076 392048
rect 517697 391990 520076 391992
rect 517697 391987 517763 391990
rect 583520 391628 584960 391868
rect 517881 391506 517947 391509
rect 517881 391504 520076 391506
rect 517881 391448 517886 391504
rect 517942 391448 520076 391504
rect 517881 391446 520076 391448
rect 517881 391443 517947 391446
rect 517697 390826 517763 390829
rect 517697 390824 520076 390826
rect 517697 390768 517702 390824
rect 517758 390768 520076 390824
rect 517697 390766 520076 390768
rect 517697 390763 517763 390766
rect 517881 390282 517947 390285
rect 517881 390280 520076 390282
rect 517881 390224 517886 390280
rect 517942 390224 520076 390280
rect 517881 390222 520076 390224
rect 517881 390219 517947 390222
rect 517697 389738 517763 389741
rect 517697 389736 520076 389738
rect 517697 389680 517702 389736
rect 517758 389680 520076 389736
rect 517697 389678 520076 389680
rect 517697 389675 517763 389678
rect 517973 389058 518039 389061
rect 517973 389056 520076 389058
rect 517973 389000 517978 389056
rect 518034 389000 520076 389056
rect 517973 388998 520076 389000
rect 517973 388995 518039 388998
rect 517881 388514 517947 388517
rect 517881 388512 520076 388514
rect 517881 388456 517886 388512
rect 517942 388456 520076 388512
rect 517881 388454 520076 388456
rect 517881 388451 517947 388454
rect 517697 387970 517763 387973
rect 517697 387968 520076 387970
rect 517697 387912 517702 387968
rect 517758 387912 520076 387968
rect 517697 387910 520076 387912
rect 517697 387907 517763 387910
rect 517881 387290 517947 387293
rect 517881 387288 520076 387290
rect 517881 387232 517886 387288
rect 517942 387232 520076 387288
rect 517881 387230 520076 387232
rect 517881 387227 517947 387230
rect 517697 386746 517763 386749
rect 517697 386744 520076 386746
rect 517697 386688 517702 386744
rect 517758 386688 520076 386744
rect 517697 386686 520076 386688
rect 517697 386683 517763 386686
rect 514017 385794 514083 385797
rect 520046 385794 520106 386172
rect 514017 385792 520106 385794
rect 514017 385736 514022 385792
rect 514078 385736 520106 385792
rect 514017 385734 520106 385736
rect 514017 385731 514083 385734
rect 451038 385188 451044 385252
rect 451108 385250 451114 385252
rect 520046 385250 520106 385492
rect 451108 385190 520106 385250
rect 451108 385188 451114 385190
rect 447726 385052 447732 385116
rect 447796 385114 447802 385116
rect 514017 385114 514083 385117
rect 447796 385112 514083 385114
rect 447796 385056 514022 385112
rect 514078 385056 514083 385112
rect 447796 385054 514083 385056
rect 447796 385052 447802 385054
rect 514017 385051 514083 385054
rect 509969 384706 510035 384709
rect 520046 384706 520106 384948
rect 509969 384704 520106 384706
rect 509969 384648 509974 384704
rect 510030 384648 520106 384704
rect 509969 384646 520106 384648
rect 509969 384643 510035 384646
rect -960 384284 480 384524
rect 449934 383964 449940 384028
rect 450004 384026 450010 384028
rect 510153 384026 510219 384029
rect 520046 384026 520106 384404
rect 450004 384024 510219 384026
rect 450004 383968 510158 384024
rect 510214 383968 510219 384024
rect 450004 383966 510219 383968
rect 450004 383964 450010 383966
rect 510153 383963 510219 383966
rect 518850 383966 520106 384026
rect 449750 383828 449756 383892
rect 449820 383890 449826 383892
rect 518850 383890 518910 383966
rect 449820 383830 518910 383890
rect 449820 383828 449826 383830
rect 447910 383692 447916 383756
rect 447980 383754 447986 383756
rect 509969 383754 510035 383757
rect 447980 383752 510035 383754
rect 447980 383696 509974 383752
rect 510030 383696 510035 383752
rect 447980 383694 510035 383696
rect 447980 383692 447986 383694
rect 509969 383691 510035 383694
rect 510153 383754 510219 383757
rect 510153 383752 520076 383754
rect 510153 383696 510158 383752
rect 510214 383696 520076 383752
rect 510153 383694 520076 383696
rect 510153 383691 510219 383694
rect 520046 382938 520106 383180
rect 509190 382878 520106 382938
rect 450854 382468 450860 382532
rect 450924 382530 450930 382532
rect 509190 382530 509250 382878
rect 518198 382604 518204 382668
rect 518268 382666 518274 382668
rect 518268 382606 520076 382666
rect 518268 382604 518274 382606
rect 450924 382470 509250 382530
rect 450924 382468 450930 382470
rect 520046 381714 520106 381956
rect 509190 381654 520106 381714
rect 448278 381108 448284 381172
rect 448348 381170 448354 381172
rect 509190 381170 509250 381654
rect 520046 381170 520106 381412
rect 448348 381110 509250 381170
rect 518850 381110 520106 381170
rect 448348 381108 448354 381110
rect 448094 380972 448100 381036
rect 448164 381034 448170 381036
rect 518850 381034 518910 381110
rect 448164 380974 518910 381034
rect 448164 380972 448170 380974
rect 518065 380898 518131 380901
rect 518065 380896 520076 380898
rect 518065 380840 518070 380896
rect 518126 380840 520076 380896
rect 518065 380838 520076 380840
rect 518065 380835 518131 380838
rect 450486 379612 450492 379676
rect 450556 379674 450562 379676
rect 520046 379674 520106 380324
rect 450556 379614 520106 379674
rect 450556 379612 450562 379614
rect 519537 379130 519603 379133
rect 550214 379130 550220 379132
rect 519537 379128 550220 379130
rect 519537 379072 519542 379128
rect 519598 379072 550220 379128
rect 519537 379070 550220 379072
rect 519537 379067 519603 379070
rect 550214 379068 550220 379070
rect 550284 379068 550290 379132
rect 517789 378994 517855 378997
rect 550398 378994 550404 378996
rect 517789 378992 550404 378994
rect 517789 378936 517794 378992
rect 517850 378936 550404 378992
rect 517789 378934 550404 378936
rect 517789 378931 517855 378934
rect 550398 378932 550404 378934
rect 550468 378932 550474 378996
rect 519721 378858 519787 378861
rect 550582 378858 550588 378860
rect 519721 378856 550588 378858
rect 519721 378800 519726 378856
rect 519782 378800 550588 378856
rect 519721 378798 550588 378800
rect 519721 378795 519787 378798
rect 550582 378796 550588 378798
rect 550652 378796 550658 378860
rect 518934 378660 518940 378724
rect 519004 378722 519010 378724
rect 550766 378722 550772 378724
rect 519004 378662 550772 378722
rect 519004 378660 519010 378662
rect 550766 378660 550772 378662
rect 550836 378660 550842 378724
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 449566 371996 449572 372060
rect 449636 372058 449642 372060
rect 518065 372058 518131 372061
rect 449636 372056 518131 372058
rect 449636 372000 518070 372056
rect 518126 372000 518131 372056
rect 449636 371998 518131 372000
rect 449636 371996 449642 371998
rect 518065 371995 518131 371998
rect 449198 371860 449204 371924
rect 449268 371922 449274 371924
rect 518198 371922 518204 371924
rect 449268 371862 518204 371922
rect 449268 371860 449274 371862
rect 518198 371860 518204 371862
rect 518268 371860 518274 371924
rect 520038 371860 520044 371924
rect 520108 371922 520114 371924
rect 564433 371922 564499 371925
rect 520108 371920 564499 371922
rect 520108 371864 564438 371920
rect 564494 371864 564499 371920
rect 520108 371862 564499 371864
rect 520108 371860 520114 371862
rect 564433 371859 564499 371862
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 223481 371242 223547 371245
rect 518014 371242 518020 371244
rect 223481 371240 518020 371242
rect 223481 371184 223486 371240
rect 223542 371184 518020 371240
rect 223481 371182 518020 371184
rect 223481 371179 223547 371182
rect 518014 371180 518020 371182
rect 518084 371180 518090 371244
rect 518525 370970 518591 370973
rect 549294 370970 549300 370972
rect 518525 370968 549300 370970
rect 518525 370912 518530 370968
rect 518586 370912 549300 370968
rect 518525 370910 549300 370912
rect 518525 370907 518591 370910
rect 549294 370908 549300 370910
rect 549364 370908 549370 370972
rect 518750 370772 518756 370836
rect 518820 370834 518826 370836
rect 550030 370834 550036 370836
rect 518820 370774 550036 370834
rect 518820 370772 518826 370774
rect 550030 370772 550036 370774
rect 550100 370772 550106 370836
rect 518341 370698 518407 370701
rect 550950 370698 550956 370700
rect 518341 370696 550956 370698
rect 518341 370640 518346 370696
rect 518402 370640 550956 370696
rect 518341 370638 550956 370640
rect 518341 370635 518407 370638
rect 550950 370636 550956 370638
rect 551020 370636 551026 370700
rect 518566 370500 518572 370564
rect 518636 370562 518642 370564
rect 553393 370562 553459 370565
rect 518636 370560 553459 370562
rect 518636 370504 553398 370560
rect 553454 370504 553459 370560
rect 518636 370502 553459 370504
rect 518636 370500 518642 370502
rect 553393 370499 553459 370502
rect 450721 369610 450787 369613
rect 450678 369608 450787 369610
rect 450678 369552 450726 369608
rect 450782 369552 450787 369608
rect 450678 369547 450787 369552
rect 450678 369036 450738 369547
rect 550081 367842 550147 367845
rect 549884 367840 550147 367842
rect 549884 367784 550086 367840
rect 550142 367784 550147 367840
rect 549884 367782 550147 367784
rect 550081 367779 550147 367782
rect 447869 367162 447935 367165
rect 447869 367160 450156 367162
rect 447869 367104 447874 367160
rect 447930 367104 450156 367160
rect 447869 367102 450156 367104
rect 447869 367099 447935 367102
rect 447869 366482 447935 366485
rect 450486 366482 450492 366484
rect 447869 366480 450492 366482
rect 447869 366424 447874 366480
rect 447930 366424 450492 366480
rect 447869 366422 450492 366424
rect 447869 366419 447935 366422
rect 450486 366420 450492 366422
rect 450556 366420 450562 366484
rect 447593 365258 447659 365261
rect 447593 365256 450156 365258
rect 447593 365200 447598 365256
rect 447654 365200 450156 365256
rect 447593 365198 450156 365200
rect 447593 365195 447659 365198
rect 580809 365122 580875 365125
rect 583520 365122 584960 365212
rect 580809 365120 584960 365122
rect 580809 365064 580814 365120
rect 580870 365064 584960 365120
rect 580809 365062 584960 365064
rect 580809 365059 580875 365062
rect 583520 364972 584960 365062
rect 549897 363898 549963 363901
rect 549854 363896 549963 363898
rect 549854 363840 549902 363896
rect 549958 363840 549963 363896
rect 549854 363835 549963 363840
rect 549854 363460 549914 363835
rect 448973 363218 449039 363221
rect 448973 363216 450156 363218
rect 448973 363160 448978 363216
rect 449034 363160 450156 363216
rect 448973 363158 450156 363160
rect 448973 363155 449039 363158
rect 449065 361314 449131 361317
rect 449065 361312 450156 361314
rect 449065 361256 449070 361312
rect 449126 361256 450156 361312
rect 449065 361254 450156 361256
rect 449065 361251 449131 361254
rect 450353 359954 450419 359957
rect 450310 359952 450419 359954
rect 450310 359896 450358 359952
rect 450414 359896 450419 359952
rect 450310 359891 450419 359896
rect 450310 359380 450370 359891
rect 551461 359138 551527 359141
rect 549884 359136 551527 359138
rect 549884 359080 551466 359136
rect 551522 359080 551527 359136
rect 549884 359078 551527 359080
rect 551461 359075 551527 359078
rect -960 358458 480 358548
rect 3049 358458 3115 358461
rect -960 358456 3115 358458
rect -960 358400 3054 358456
rect 3110 358400 3115 358456
rect -960 358398 3115 358400
rect -960 358308 480 358398
rect 3049 358395 3115 358398
rect 450261 357642 450327 357645
rect 450261 357640 450370 357642
rect 450261 357584 450266 357640
rect 450322 357584 450370 357640
rect 450261 357579 450370 357584
rect 450310 357340 450370 357579
rect 447685 355466 447751 355469
rect 447685 355464 450156 355466
rect 447685 355408 447690 355464
rect 447746 355408 450156 355464
rect 447685 355406 450156 355408
rect 447685 355403 447751 355406
rect 551369 354786 551435 354789
rect 549884 354784 551435 354786
rect 549884 354728 551374 354784
rect 551430 354728 551435 354784
rect 549884 354726 551435 354728
rect 551369 354723 551435 354726
rect 450169 354106 450235 354109
rect 450126 354104 450235 354106
rect 450126 354048 450174 354104
rect 450230 354048 450235 354104
rect 450126 354043 450235 354048
rect 450126 353532 450186 354043
rect 450077 351930 450143 351933
rect 579613 351930 579679 351933
rect 583520 351930 584960 352020
rect 450077 351928 450186 351930
rect 450077 351872 450082 351928
rect 450138 351872 450186 351928
rect 450077 351867 450186 351872
rect 579613 351928 584960 351930
rect 579613 351872 579618 351928
rect 579674 351872 584960 351928
rect 579613 351870 584960 351872
rect 579613 351867 579679 351870
rect 450126 351492 450186 351867
rect 583520 351780 584960 351870
rect 550081 350434 550147 350437
rect 549884 350432 550147 350434
rect 549884 350376 550086 350432
rect 550142 350376 550147 350432
rect 549884 350374 550147 350376
rect 550081 350371 550147 350374
rect 449985 350162 450051 350165
rect 449985 350160 450186 350162
rect 449985 350104 449990 350160
rect 450046 350104 450186 350160
rect 449985 350102 450186 350104
rect 449985 350099 450051 350102
rect 450126 349588 450186 350102
rect 449893 347850 449959 347853
rect 449893 347848 450186 347850
rect 449893 347792 449898 347848
rect 449954 347792 450186 347848
rect 449893 347790 450186 347792
rect 449893 347787 449959 347790
rect 450126 347684 450186 347790
rect 551277 345946 551343 345949
rect 549884 345944 551343 345946
rect 549884 345888 551282 345944
rect 551338 345888 551343 345944
rect 549884 345886 551343 345888
rect 551277 345883 551343 345886
rect 447777 345810 447843 345813
rect 447777 345808 450156 345810
rect 447777 345752 447782 345808
rect 447838 345752 450156 345808
rect 447777 345750 450156 345752
rect 447777 345747 447843 345750
rect -960 345402 480 345492
rect 2957 345402 3023 345405
rect -960 345400 3023 345402
rect -960 345344 2962 345400
rect 3018 345344 3023 345400
rect -960 345342 3023 345344
rect -960 345252 480 345342
rect 2957 345339 3023 345342
rect 449157 343770 449223 343773
rect 449157 343768 450156 343770
rect 449157 343712 449162 343768
rect 449218 343712 450156 343768
rect 449157 343710 450156 343712
rect 449157 343707 449223 343710
rect 449341 341866 449407 341869
rect 449341 341864 450156 341866
rect 449341 341808 449346 341864
rect 449402 341808 450156 341864
rect 449341 341806 450156 341808
rect 449341 341803 449407 341806
rect 552473 341594 552539 341597
rect 549884 341592 552539 341594
rect 549884 341536 552478 341592
rect 552534 341536 552539 341592
rect 549884 341534 552539 341536
rect 552473 341531 552539 341534
rect 449249 339962 449315 339965
rect 449249 339960 450156 339962
rect 449249 339904 449254 339960
rect 449310 339904 450156 339960
rect 449249 339902 450156 339904
rect 449249 339899 449315 339902
rect 583520 338452 584960 338692
rect 449525 337922 449591 337925
rect 449525 337920 450156 337922
rect 449525 337864 449530 337920
rect 449586 337864 450156 337920
rect 449525 337862 450156 337864
rect 449525 337859 449591 337862
rect 552381 337242 552447 337245
rect 549884 337240 552447 337242
rect 549884 337184 552386 337240
rect 552442 337184 552447 337240
rect 549884 337182 552447 337184
rect 552381 337179 552447 337182
rect 449617 336018 449683 336021
rect 449617 336016 450156 336018
rect 449617 335960 449622 336016
rect 449678 335960 450156 336016
rect 449617 335958 450156 335960
rect 449617 335955 449683 335958
rect 449433 334114 449499 334117
rect 449433 334112 450156 334114
rect 449433 334056 449438 334112
rect 449494 334056 450156 334112
rect 449433 334054 450156 334056
rect 449433 334051 449499 334054
rect 552289 332890 552355 332893
rect 549884 332888 552355 332890
rect 549884 332832 552294 332888
rect 552350 332832 552355 332888
rect 549884 332830 552355 332832
rect 552289 332827 552355 332830
rect -960 332196 480 332436
rect 449709 332074 449775 332077
rect 449709 332072 450156 332074
rect 449709 332016 449714 332072
rect 449770 332016 450156 332072
rect 449709 332014 450156 332016
rect 449709 332011 449775 332014
rect 449801 330170 449867 330173
rect 449801 330168 450156 330170
rect 449801 330112 449806 330168
rect 449862 330112 450156 330168
rect 449801 330110 450156 330112
rect 449801 330107 449867 330110
rect 552197 328538 552263 328541
rect 549884 328536 552263 328538
rect 549884 328480 552202 328536
rect 552258 328480 552263 328536
rect 549884 328478 552263 328480
rect 552197 328475 552263 328478
rect 449382 328204 449388 328268
rect 449452 328266 449458 328268
rect 449452 328206 450156 328266
rect 449452 328204 449458 328206
rect 447961 326226 448027 326229
rect 447961 326224 450156 326226
rect 447961 326168 447966 326224
rect 448022 326168 450156 326224
rect 447961 326166 450156 326168
rect 447961 326163 448027 326166
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 448145 324322 448211 324325
rect 448145 324320 450156 324322
rect 448145 324264 448150 324320
rect 448206 324264 450156 324320
rect 448145 324262 450156 324264
rect 448145 324259 448211 324262
rect 552105 324050 552171 324053
rect 549884 324048 552171 324050
rect 549884 323992 552110 324048
rect 552166 323992 552171 324048
rect 549884 323990 552171 323992
rect 552105 323987 552171 323990
rect 448053 322418 448119 322421
rect 448053 322416 450156 322418
rect 448053 322360 448058 322416
rect 448114 322360 450156 322416
rect 448053 322358 450156 322360
rect 448053 322355 448119 322358
rect 448237 320514 448303 320517
rect 448237 320512 450156 320514
rect 448237 320456 448242 320512
rect 448298 320456 450156 320512
rect 448237 320454 450156 320456
rect 448237 320451 448303 320454
rect 552013 319698 552079 319701
rect 549884 319696 552079 319698
rect 549884 319640 552018 319696
rect 552074 319640 552079 319696
rect 549884 319638 552079 319640
rect 552013 319635 552079 319638
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 448329 318474 448395 318477
rect 448329 318472 450156 318474
rect 448329 318416 448334 318472
rect 448390 318416 450156 318472
rect 448329 318414 450156 318416
rect 448329 318411 448395 318414
rect 448421 316570 448487 316573
rect 448421 316568 450156 316570
rect 448421 316512 448426 316568
rect 448482 316512 450156 316568
rect 448421 316510 450156 316512
rect 448421 316507 448487 316510
rect 549345 315754 549411 315757
rect 549302 315752 549411 315754
rect 549302 315696 549350 315752
rect 549406 315696 549411 315752
rect 549302 315691 549411 315696
rect 549302 315316 549362 315691
rect 447726 314604 447732 314668
rect 447796 314666 447802 314668
rect 447796 314606 450156 314666
rect 447796 314604 447802 314606
rect 447910 312564 447916 312628
rect 447980 312626 447986 312628
rect 447980 312566 450156 312626
rect 447980 312564 447986 312566
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 449934 311204 449940 311268
rect 450004 311266 450010 311268
rect 450004 311206 450186 311266
rect 450004 311204 450010 311206
rect 450126 310692 450186 311206
rect 551185 310994 551251 310997
rect 549884 310992 551251 310994
rect 549884 310936 551190 310992
rect 551246 310936 551251 310992
rect 549884 310934 551251 310936
rect 551185 310931 551251 310934
rect 449198 308756 449204 308820
rect 449268 308818 449274 308820
rect 449268 308758 450156 308818
rect 449268 308756 449274 308758
rect 549345 307186 549411 307189
rect 549302 307184 549411 307186
rect 549302 307128 549350 307184
rect 549406 307128 549411 307184
rect 549302 307123 549411 307128
rect 448094 306716 448100 306780
rect 448164 306778 448170 306780
rect 448164 306718 450156 306778
rect 448164 306716 448170 306718
rect 549302 306612 549362 307123
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 448278 304812 448284 304876
rect 448348 304874 448354 304876
rect 448348 304814 450156 304874
rect 448348 304812 448354 304814
rect 447777 302970 447843 302973
rect 449566 302970 449572 302972
rect 447777 302968 449572 302970
rect 447777 302912 447782 302968
rect 447838 302912 449572 302968
rect 447777 302910 449572 302912
rect 447777 302907 447843 302910
rect 449566 302908 449572 302910
rect 449636 302970 449642 302972
rect 449636 302910 450156 302970
rect 449636 302908 449642 302910
rect 551093 302290 551159 302293
rect 549884 302288 551159 302290
rect 549884 302232 551098 302288
rect 551154 302232 551159 302288
rect 549884 302230 551159 302232
rect 551093 302227 551159 302230
rect 447869 301066 447935 301069
rect 447869 301064 450156 301066
rect 447869 301008 447874 301064
rect 447930 301008 450156 301064
rect 447869 301006 450156 301008
rect 447869 301003 447935 301006
rect 450854 299508 450860 299572
rect 450924 299570 450930 299572
rect 451457 299570 451523 299573
rect 450924 299568 451523 299570
rect 450924 299512 451462 299568
rect 451518 299512 451523 299568
rect 450924 299510 451523 299512
rect 450924 299508 450930 299510
rect 451457 299507 451523 299510
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 548609 298074 548675 298077
rect 553761 298074 553827 298077
rect 548609 298072 553827 298074
rect 548609 298016 548614 298072
rect 548670 298016 553766 298072
rect 553822 298016 553827 298072
rect 548609 298014 553827 298016
rect 548609 298011 548675 298014
rect 553761 298011 553827 298014
rect 449750 297876 449756 297940
rect 449820 297938 449826 297940
rect 454493 297938 454559 297941
rect 449820 297936 454559 297938
rect 449820 297880 454498 297936
rect 454554 297880 454559 297936
rect 449820 297878 454559 297880
rect 449820 297876 449826 297878
rect 454493 297875 454559 297878
rect 488901 297938 488967 297941
rect 550766 297938 550772 297940
rect 488901 297936 550772 297938
rect 488901 297880 488906 297936
rect 488962 297880 550772 297936
rect 488901 297878 550772 297880
rect 488901 297875 488967 297878
rect 550766 297876 550772 297878
rect 550836 297876 550842 297940
rect 451038 297740 451044 297804
rect 451108 297802 451114 297804
rect 457621 297802 457687 297805
rect 451108 297800 457687 297802
rect 451108 297744 457626 297800
rect 457682 297744 457687 297800
rect 451108 297742 457687 297744
rect 451108 297740 451114 297742
rect 457621 297739 457687 297742
rect 492029 297802 492095 297805
rect 550582 297802 550588 297804
rect 492029 297800 550588 297802
rect 492029 297744 492034 297800
rect 492090 297744 550588 297800
rect 492029 297742 550588 297744
rect 492029 297739 492095 297742
rect 550582 297740 550588 297742
rect 550652 297740 550658 297804
rect 495157 297666 495223 297669
rect 550214 297666 550220 297668
rect 495157 297664 550220 297666
rect 495157 297608 495162 297664
rect 495218 297608 550220 297664
rect 495157 297606 550220 297608
rect 495157 297603 495223 297606
rect 550214 297604 550220 297606
rect 550284 297604 550290 297668
rect 532693 297530 532759 297533
rect 548926 297530 548932 297532
rect 532693 297528 548932 297530
rect 532693 297472 532698 297528
rect 532754 297472 548932 297528
rect 532693 297470 548932 297472
rect 532693 297467 532759 297470
rect 548926 297468 548932 297470
rect 548996 297468 549002 297532
rect 529565 297394 529631 297397
rect 550950 297394 550956 297396
rect 529565 297392 550956 297394
rect 529565 297336 529570 297392
rect 529626 297336 550956 297392
rect 529565 297334 550956 297336
rect 529565 297331 529631 297334
rect 550950 297332 550956 297334
rect 551020 297332 551026 297396
rect 485773 297258 485839 297261
rect 550398 297258 550404 297260
rect 485773 297256 550404 297258
rect 485773 297200 485778 297256
rect 485834 297200 550404 297256
rect 485773 297198 550404 297200
rect 485773 297195 485839 297198
rect 550398 297196 550404 297198
rect 550468 297196 550474 297260
rect -960 293178 480 293268
rect 3233 293178 3299 293181
rect -960 293176 3299 293178
rect -960 293120 3238 293176
rect 3294 293120 3299 293176
rect -960 293118 3299 293120
rect -960 293028 480 293118
rect 3233 293115 3299 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3325 267202 3391 267205
rect -960 267200 3391 267202
rect -960 267144 3330 267200
rect 3386 267144 3391 267200
rect -960 267142 3391 267144
rect -960 267052 480 267142
rect 3325 267139 3391 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 2957 254146 3023 254149
rect -960 254144 3023 254146
rect -960 254088 2962 254144
rect 3018 254088 3023 254144
rect -960 254086 3023 254088
rect -960 253996 480 254086
rect 2957 254083 3023 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3785 241090 3851 241093
rect -960 241088 3851 241090
rect -960 241032 3790 241088
rect 3846 241032 3851 241088
rect -960 241030 3851 241032
rect -960 240940 480 241030
rect 3785 241027 3851 241030
rect 580717 232386 580783 232389
rect 583520 232386 584960 232476
rect 580717 232384 584960 232386
rect 580717 232328 580722 232384
rect 580778 232328 584960 232384
rect 580717 232326 584960 232328
rect 580717 232323 580783 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580625 219058 580691 219061
rect 583520 219058 584960 219148
rect 580625 219056 584960 219058
rect 580625 219000 580630 219056
rect 580686 219000 584960 219056
rect 580625 218998 584960 219000
rect 580625 218995 580691 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3693 201922 3759 201925
rect -960 201920 3759 201922
rect -960 201864 3698 201920
rect 3754 201864 3759 201920
rect -960 201862 3759 201864
rect -960 201772 480 201862
rect 3693 201859 3759 201862
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 579613 179210 579679 179213
rect 583520 179210 584960 179300
rect 579613 179208 584960 179210
rect 579613 179152 579618 179208
rect 579674 179152 584960 179208
rect 579613 179150 584960 179152
rect 579613 179147 579679 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect 580533 152690 580599 152693
rect 583520 152690 584960 152780
rect 580533 152688 584960 152690
rect 580533 152632 580538 152688
rect 580594 152632 584960 152688
rect 580533 152630 584960 152632
rect 580533 152627 580599 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 580441 139362 580507 139365
rect 583520 139362 584960 139452
rect 580441 139360 584960 139362
rect 580441 139304 580446 139360
rect 580502 139304 584960 139360
rect 580441 139302 584960 139304
rect 580441 139299 580507 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579613 112842 579679 112845
rect 583520 112842 584960 112932
rect 579613 112840 584960 112842
rect 579613 112784 579618 112840
rect 579674 112784 584960 112840
rect 579613 112782 584960 112784
rect 579613 112779 579679 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3877 110666 3943 110669
rect -960 110664 3943 110666
rect -960 110608 3882 110664
rect 3938 110608 3943 110664
rect -960 110606 3943 110608
rect -960 110516 480 110606
rect 3877 110603 3943 110606
rect 580349 99514 580415 99517
rect 583520 99514 584960 99604
rect 580349 99512 584960 99514
rect 580349 99456 580354 99512
rect 580410 99456 584960 99512
rect 580349 99454 584960 99456
rect 580349 99451 580415 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2957 84690 3023 84693
rect -960 84688 3023 84690
rect -960 84632 2962 84688
rect 3018 84632 3023 84688
rect -960 84630 3023 84632
rect -960 84540 480 84630
rect 2957 84627 3023 84630
rect 169753 79930 169819 79933
rect 170259 79930 170325 79933
rect 169753 79928 170325 79930
rect 169753 79872 169758 79928
rect 169814 79872 170264 79928
rect 170320 79872 170325 79928
rect 169753 79870 170325 79872
rect 169753 79867 169819 79870
rect 170259 79867 170325 79870
rect 142153 77482 142219 77485
rect 142521 77482 142587 77485
rect 142153 77480 142587 77482
rect 142153 77424 142158 77480
rect 142214 77424 142526 77480
rect 142582 77424 142587 77480
rect 142153 77422 142587 77424
rect 142153 77419 142219 77422
rect 142521 77419 142587 77422
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3693 71634 3759 71637
rect -960 71632 3759 71634
rect -960 71576 3698 71632
rect 3754 71576 3759 71632
rect -960 71574 3759 71576
rect -960 71484 480 71574
rect 3693 71571 3759 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 550081 46884 550147 46885
rect 550030 46882 550036 46884
rect 549990 46822 550036 46882
rect 550100 46880 550147 46884
rect 550142 46824 550147 46880
rect 550030 46820 550036 46822
rect 550100 46820 550147 46824
rect 550081 46819 550147 46820
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3785 32466 3851 32469
rect -960 32464 3851 32466
rect -960 32408 3790 32464
rect 3846 32408 3851 32464
rect -960 32406 3851 32408
rect -960 32316 480 32406
rect 3785 32403 3851 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect -960 6430 674 6490
rect 583520 6476 584960 6566
rect -960 6354 480 6430
rect 614 6354 674 6430
rect -960 6340 674 6354
rect 246 6294 674 6340
rect 246 5810 306 6294
rect 246 5750 6930 5810
rect 6870 5674 6930 5750
rect 558862 5674 558868 5676
rect 6870 5614 558868 5674
rect 558862 5612 558868 5614
rect 558932 5612 558938 5676
<< via3 >>
rect 518020 422996 518084 423060
rect 518756 420412 518820 420476
rect 558868 419868 558932 419932
rect 519860 419384 519924 419388
rect 519860 419328 519910 419384
rect 519910 419328 519924 419384
rect 519860 419324 519924 419328
rect 518572 418508 518636 418572
rect 518940 397292 519004 397356
rect 449388 393484 449452 393548
rect 451044 385188 451108 385252
rect 447732 385052 447796 385116
rect 449940 383964 450004 384028
rect 449756 383828 449820 383892
rect 447916 383692 447980 383756
rect 450860 382468 450924 382532
rect 518204 382604 518268 382668
rect 448284 381108 448348 381172
rect 448100 380972 448164 381036
rect 450492 379612 450556 379676
rect 550220 379068 550284 379132
rect 550404 378932 550468 378996
rect 550588 378796 550652 378860
rect 518940 378660 519004 378724
rect 550772 378660 550836 378724
rect 449572 371996 449636 372060
rect 449204 371860 449268 371924
rect 518204 371860 518268 371924
rect 520044 371860 520108 371924
rect 518020 371180 518084 371244
rect 549300 370908 549364 370972
rect 518756 370772 518820 370836
rect 550036 370772 550100 370836
rect 550956 370636 551020 370700
rect 518572 370500 518636 370564
rect 450492 366420 450556 366484
rect 449388 328204 449452 328268
rect 447732 314604 447796 314668
rect 447916 312564 447980 312628
rect 449940 311204 450004 311268
rect 449204 308756 449268 308820
rect 448100 306716 448164 306780
rect 448284 304812 448348 304876
rect 449572 302908 449636 302972
rect 450860 299508 450924 299572
rect 449756 297876 449820 297940
rect 550772 297876 550836 297940
rect 451044 297740 451108 297804
rect 550588 297740 550652 297804
rect 550220 297604 550284 297668
rect 548932 297468 548996 297532
rect 550956 297332 551020 297396
rect 550404 297196 550468 297260
rect 550036 46880 550100 46884
rect 550036 46824 550086 46880
rect 550086 46824 550100 46880
rect 550036 46820 550100 46824
rect 558868 5612 558932 5676
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 202000 78134 222618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 202000 81854 226338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 202000 85574 230058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 202000 92414 236898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 202000 96134 204618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 202000 99854 208338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 202000 103574 212058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 202000 110414 218898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 202000 114134 222618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 202000 117854 226338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 202000 121574 230058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 202000 128414 236898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 202000 132134 204618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 202000 135854 208338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 202000 139574 212058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 202000 146414 218898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 202000 150134 222618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 202000 153854 226338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 202000 157574 230058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 202000 164414 236898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 202000 168134 204618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 202000 171854 208338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 202000 175574 212058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 202000 182414 218898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 202000 186134 222618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 202000 189854 226338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 202000 193574 230058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 202000 200414 236898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 202000 204134 204618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 202000 207854 208338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 202000 211574 212058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 202000 218414 218898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 202000 222134 222618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 202000 225854 226338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 202000 229574 230058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 202000 236414 236898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 202000 240134 204618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 202000 243854 208338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 202000 247574 212058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 202000 254414 218898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 202000 258134 222618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 202000 261854 226338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 84208 183454 84528 183486
rect 84208 183218 84250 183454
rect 84486 183218 84528 183454
rect 84208 183134 84528 183218
rect 84208 182898 84250 183134
rect 84486 182898 84528 183134
rect 84208 182866 84528 182898
rect 114928 183454 115248 183486
rect 114928 183218 114970 183454
rect 115206 183218 115248 183454
rect 114928 183134 115248 183218
rect 114928 182898 114970 183134
rect 115206 182898 115248 183134
rect 114928 182866 115248 182898
rect 145648 183454 145968 183486
rect 145648 183218 145690 183454
rect 145926 183218 145968 183454
rect 145648 183134 145968 183218
rect 145648 182898 145690 183134
rect 145926 182898 145968 183134
rect 145648 182866 145968 182898
rect 176368 183454 176688 183486
rect 176368 183218 176410 183454
rect 176646 183218 176688 183454
rect 176368 183134 176688 183218
rect 176368 182898 176410 183134
rect 176646 182898 176688 183134
rect 176368 182866 176688 182898
rect 207088 183454 207408 183486
rect 207088 183218 207130 183454
rect 207366 183218 207408 183454
rect 207088 183134 207408 183218
rect 207088 182898 207130 183134
rect 207366 182898 207408 183134
rect 207088 182866 207408 182898
rect 237808 183454 238128 183486
rect 237808 183218 237850 183454
rect 238086 183218 238128 183454
rect 237808 183134 238128 183218
rect 237808 182898 237850 183134
rect 238086 182898 238128 183134
rect 237808 182866 238128 182898
rect 99568 165454 99888 165486
rect 99568 165218 99610 165454
rect 99846 165218 99888 165454
rect 99568 165134 99888 165218
rect 99568 164898 99610 165134
rect 99846 164898 99888 165134
rect 99568 164866 99888 164898
rect 130288 165454 130608 165486
rect 130288 165218 130330 165454
rect 130566 165218 130608 165454
rect 130288 165134 130608 165218
rect 130288 164898 130330 165134
rect 130566 164898 130608 165134
rect 130288 164866 130608 164898
rect 161008 165454 161328 165486
rect 161008 165218 161050 165454
rect 161286 165218 161328 165454
rect 161008 165134 161328 165218
rect 161008 164898 161050 165134
rect 161286 164898 161328 165134
rect 161008 164866 161328 164898
rect 191728 165454 192048 165486
rect 191728 165218 191770 165454
rect 192006 165218 192048 165454
rect 191728 165134 192048 165218
rect 191728 164898 191770 165134
rect 192006 164898 192048 165134
rect 191728 164866 192048 164898
rect 222448 165454 222768 165486
rect 222448 165218 222490 165454
rect 222726 165218 222768 165454
rect 222448 165134 222768 165218
rect 222448 164898 222490 165134
rect 222726 164898 222768 165134
rect 222448 164866 222768 164898
rect 253168 165454 253488 165486
rect 253168 165218 253210 165454
rect 253446 165218 253488 165454
rect 253168 165134 253488 165218
rect 253168 164898 253210 165134
rect 253446 164898 253488 165134
rect 253168 164866 253488 164898
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 84208 147454 84528 147486
rect 84208 147218 84250 147454
rect 84486 147218 84528 147454
rect 84208 147134 84528 147218
rect 84208 146898 84250 147134
rect 84486 146898 84528 147134
rect 84208 146866 84528 146898
rect 114928 147454 115248 147486
rect 114928 147218 114970 147454
rect 115206 147218 115248 147454
rect 114928 147134 115248 147218
rect 114928 146898 114970 147134
rect 115206 146898 115248 147134
rect 114928 146866 115248 146898
rect 145648 147454 145968 147486
rect 145648 147218 145690 147454
rect 145926 147218 145968 147454
rect 145648 147134 145968 147218
rect 145648 146898 145690 147134
rect 145926 146898 145968 147134
rect 145648 146866 145968 146898
rect 176368 147454 176688 147486
rect 176368 147218 176410 147454
rect 176646 147218 176688 147454
rect 176368 147134 176688 147218
rect 176368 146898 176410 147134
rect 176646 146898 176688 147134
rect 176368 146866 176688 146898
rect 207088 147454 207408 147486
rect 207088 147218 207130 147454
rect 207366 147218 207408 147454
rect 207088 147134 207408 147218
rect 207088 146898 207130 147134
rect 207366 146898 207408 147134
rect 207088 146866 207408 146898
rect 237808 147454 238128 147486
rect 237808 147218 237850 147454
rect 238086 147218 238128 147454
rect 237808 147134 238128 147218
rect 237808 146898 237850 147134
rect 238086 146898 238128 147134
rect 237808 146866 238128 146898
rect 99568 129454 99888 129486
rect 99568 129218 99610 129454
rect 99846 129218 99888 129454
rect 99568 129134 99888 129218
rect 99568 128898 99610 129134
rect 99846 128898 99888 129134
rect 99568 128866 99888 128898
rect 130288 129454 130608 129486
rect 130288 129218 130330 129454
rect 130566 129218 130608 129454
rect 130288 129134 130608 129218
rect 130288 128898 130330 129134
rect 130566 128898 130608 129134
rect 130288 128866 130608 128898
rect 161008 129454 161328 129486
rect 161008 129218 161050 129454
rect 161286 129218 161328 129454
rect 161008 129134 161328 129218
rect 161008 128898 161050 129134
rect 161286 128898 161328 129134
rect 161008 128866 161328 128898
rect 191728 129454 192048 129486
rect 191728 129218 191770 129454
rect 192006 129218 192048 129454
rect 191728 129134 192048 129218
rect 191728 128898 191770 129134
rect 192006 128898 192048 129134
rect 191728 128866 192048 128898
rect 222448 129454 222768 129486
rect 222448 129218 222490 129454
rect 222726 129218 222768 129454
rect 222448 129134 222768 129218
rect 222448 128898 222490 129134
rect 222726 128898 222768 129134
rect 222448 128866 222768 128898
rect 253168 129454 253488 129486
rect 253168 129218 253210 129454
rect 253446 129218 253488 129454
rect 253168 129134 253488 129218
rect 253168 128898 253210 129134
rect 253446 128898 253488 129134
rect 253168 128866 253488 128898
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 84208 111454 84528 111486
rect 84208 111218 84250 111454
rect 84486 111218 84528 111454
rect 84208 111134 84528 111218
rect 84208 110898 84250 111134
rect 84486 110898 84528 111134
rect 84208 110866 84528 110898
rect 114928 111454 115248 111486
rect 114928 111218 114970 111454
rect 115206 111218 115248 111454
rect 114928 111134 115248 111218
rect 114928 110898 114970 111134
rect 115206 110898 115248 111134
rect 114928 110866 115248 110898
rect 145648 111454 145968 111486
rect 145648 111218 145690 111454
rect 145926 111218 145968 111454
rect 145648 111134 145968 111218
rect 145648 110898 145690 111134
rect 145926 110898 145968 111134
rect 145648 110866 145968 110898
rect 176368 111454 176688 111486
rect 176368 111218 176410 111454
rect 176646 111218 176688 111454
rect 176368 111134 176688 111218
rect 176368 110898 176410 111134
rect 176646 110898 176688 111134
rect 176368 110866 176688 110898
rect 207088 111454 207408 111486
rect 207088 111218 207130 111454
rect 207366 111218 207408 111454
rect 207088 111134 207408 111218
rect 207088 110898 207130 111134
rect 207366 110898 207408 111134
rect 207088 110866 207408 110898
rect 237808 111454 238128 111486
rect 237808 111218 237850 111454
rect 238086 111218 238128 111454
rect 237808 111134 238128 111218
rect 237808 110898 237850 111134
rect 238086 110898 238128 111134
rect 237808 110866 238128 110898
rect 99568 93454 99888 93486
rect 99568 93218 99610 93454
rect 99846 93218 99888 93454
rect 99568 93134 99888 93218
rect 99568 92898 99610 93134
rect 99846 92898 99888 93134
rect 99568 92866 99888 92898
rect 130288 93454 130608 93486
rect 130288 93218 130330 93454
rect 130566 93218 130608 93454
rect 130288 93134 130608 93218
rect 130288 92898 130330 93134
rect 130566 92898 130608 93134
rect 130288 92866 130608 92898
rect 161008 93454 161328 93486
rect 161008 93218 161050 93454
rect 161286 93218 161328 93454
rect 161008 93134 161328 93218
rect 161008 92898 161050 93134
rect 161286 92898 161328 93134
rect 161008 92866 161328 92898
rect 191728 93454 192048 93486
rect 191728 93218 191770 93454
rect 192006 93218 192048 93454
rect 191728 93134 192048 93218
rect 191728 92898 191770 93134
rect 192006 92898 192048 93134
rect 191728 92866 192048 92898
rect 222448 93454 222768 93486
rect 222448 93218 222490 93454
rect 222726 93218 222768 93454
rect 222448 93134 222768 93218
rect 222448 92898 222490 93134
rect 222726 92898 222768 93134
rect 222448 92866 222768 92898
rect 253168 93454 253488 93486
rect 253168 93218 253210 93454
rect 253446 93218 253488 93454
rect 253168 93134 253488 93218
rect 253168 92898 253210 93134
rect 253446 92898 253488 93134
rect 253168 92866 253488 92898
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 78000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 78000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 78000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 78000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 78000
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 78000
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 78000
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 78000
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 78000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 78000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 78000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 78000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 78000
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 78000
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 78000
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 78000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 78000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 78000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 78000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 78000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 78000
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 78000
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 68614 175574 78000
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 78000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 78000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 78000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 78000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 61174 204134 78000
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 78000
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 78000
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 78000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 78000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 78000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 78000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 78000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 78000
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 78000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 78000
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 75454 254414 78000
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 78000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 78000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 449387 393548 449453 393549
rect 449387 393484 449388 393548
rect 449452 393484 449453 393548
rect 449387 393483 449453 393484
rect 447731 385116 447797 385117
rect 447731 385052 447732 385116
rect 447796 385052 447797 385116
rect 447731 385051 447797 385052
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 447734 314669 447794 385051
rect 447915 383756 447981 383757
rect 447915 383692 447916 383756
rect 447980 383692 447981 383756
rect 447915 383691 447981 383692
rect 447731 314668 447797 314669
rect 447731 314604 447732 314668
rect 447796 314604 447797 314668
rect 447731 314603 447797 314604
rect 447918 312629 447978 383691
rect 448283 381172 448349 381173
rect 448283 381108 448284 381172
rect 448348 381108 448349 381172
rect 448283 381107 448349 381108
rect 448099 381036 448165 381037
rect 448099 380972 448100 381036
rect 448164 380972 448165 381036
rect 448099 380971 448165 380972
rect 447915 312628 447981 312629
rect 447915 312564 447916 312628
rect 447980 312564 447981 312628
rect 447915 312563 447981 312564
rect 448102 306781 448162 380971
rect 448099 306780 448165 306781
rect 448099 306716 448100 306780
rect 448164 306716 448165 306780
rect 448099 306715 448165 306716
rect 448286 304877 448346 381107
rect 449203 371924 449269 371925
rect 449203 371860 449204 371924
rect 449268 371860 449269 371924
rect 449203 371859 449269 371860
rect 449206 308821 449266 371859
rect 449390 328269 449450 393483
rect 451043 385252 451109 385253
rect 451043 385188 451044 385252
rect 451108 385188 451109 385252
rect 451043 385187 451109 385188
rect 449939 384028 450005 384029
rect 449939 383964 449940 384028
rect 450004 383964 450005 384028
rect 449939 383963 450005 383964
rect 449755 383892 449821 383893
rect 449755 383828 449756 383892
rect 449820 383828 449821 383892
rect 449755 383827 449821 383828
rect 449571 372060 449637 372061
rect 449571 371996 449572 372060
rect 449636 371996 449637 372060
rect 449571 371995 449637 371996
rect 449387 328268 449453 328269
rect 449387 328204 449388 328268
rect 449452 328204 449453 328268
rect 449387 328203 449453 328204
rect 449203 308820 449269 308821
rect 449203 308756 449204 308820
rect 449268 308756 449269 308820
rect 449203 308755 449269 308756
rect 448283 304876 448349 304877
rect 448283 304812 448284 304876
rect 448348 304812 448349 304876
rect 448283 304811 448349 304812
rect 449574 302973 449634 371995
rect 449571 302972 449637 302973
rect 449571 302908 449572 302972
rect 449636 302908 449637 302972
rect 449571 302907 449637 302908
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 449758 297941 449818 383827
rect 449942 311269 450002 383963
rect 450859 382532 450925 382533
rect 450859 382468 450860 382532
rect 450924 382468 450925 382532
rect 450859 382467 450925 382468
rect 450491 379676 450557 379677
rect 450491 379612 450492 379676
rect 450556 379612 450557 379676
rect 450491 379611 450557 379612
rect 450494 366485 450554 379611
rect 450491 366484 450557 366485
rect 450491 366420 450492 366484
rect 450556 366420 450557 366484
rect 450491 366419 450557 366420
rect 449939 311268 450005 311269
rect 449939 311204 449940 311268
rect 450004 311204 450005 311268
rect 449939 311203 450005 311204
rect 450862 299573 450922 382467
rect 450859 299572 450925 299573
rect 450859 299508 450860 299572
rect 450924 299508 450925 299572
rect 450859 299507 450925 299508
rect 449755 297940 449821 297941
rect 449755 297876 449756 297940
rect 449820 297876 449821 297940
rect 449755 297875 449821 297876
rect 451046 297805 451106 385187
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 372000 452414 380898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 372000 456134 384618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 372000 459854 388338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 372000 463574 392058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 372000 470414 398898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 372000 474134 402618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 372000 477854 406338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 372000 481574 374058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 372000 488414 380898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 372000 492134 384618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 372000 495854 388338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 372000 499574 392058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 372000 506414 398898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 372000 510134 402618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 372000 513854 406338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 518019 423060 518085 423061
rect 518019 422996 518020 423060
rect 518084 422996 518085 423060
rect 518019 422995 518085 422996
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 372000 517574 374058
rect 518022 371245 518082 422995
rect 523794 422000 524414 452898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 422000 528134 456618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 422000 531854 424338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 422000 535574 428058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 422000 542414 434898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 422000 546134 438618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 422000 549854 442338
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 422000 553574 446058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 422000 560414 452898
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 518755 420476 518821 420477
rect 518755 420412 518756 420476
rect 518820 420412 518821 420476
rect 518755 420411 518821 420412
rect 518571 418572 518637 418573
rect 518571 418508 518572 418572
rect 518636 418508 518637 418572
rect 518571 418507 518637 418508
rect 518203 382668 518269 382669
rect 518203 382604 518204 382668
rect 518268 382604 518269 382668
rect 518203 382603 518269 382604
rect 518206 371925 518266 382603
rect 518203 371924 518269 371925
rect 518203 371860 518204 371924
rect 518268 371860 518269 371924
rect 518203 371859 518269 371860
rect 518019 371244 518085 371245
rect 518019 371180 518020 371244
rect 518084 371180 518085 371244
rect 518019 371179 518085 371180
rect 518574 370565 518634 418507
rect 518758 370837 518818 420411
rect 558867 419932 558933 419933
rect 558867 419868 558868 419932
rect 558932 419868 558933 419932
rect 558867 419867 558933 419868
rect 519859 419388 519925 419389
rect 519859 419324 519860 419388
rect 519924 419324 519925 419388
rect 519859 419323 519925 419324
rect 519862 412650 519922 419323
rect 539568 417454 539888 417486
rect 539568 417218 539610 417454
rect 539846 417218 539888 417454
rect 539568 417134 539888 417218
rect 539568 416898 539610 417134
rect 539846 416898 539888 417134
rect 539568 416866 539888 416898
rect 519862 412590 520106 412650
rect 518939 397356 519005 397357
rect 518939 397292 518940 397356
rect 519004 397292 519005 397356
rect 518939 397291 519005 397292
rect 518942 378725 519002 397291
rect 518939 378724 519005 378725
rect 518939 378660 518940 378724
rect 519004 378660 519005 378724
rect 518939 378659 519005 378660
rect 520046 371925 520106 412590
rect 524208 399454 524528 399486
rect 524208 399218 524250 399454
rect 524486 399218 524528 399454
rect 524208 399134 524528 399218
rect 524208 398898 524250 399134
rect 524486 398898 524528 399134
rect 524208 398866 524528 398898
rect 554928 399454 555248 399486
rect 554928 399218 554970 399454
rect 555206 399218 555248 399454
rect 554928 399134 555248 399218
rect 554928 398898 554970 399134
rect 555206 398898 555248 399134
rect 554928 398866 555248 398898
rect 550219 379132 550285 379133
rect 550219 379068 550220 379132
rect 550284 379068 550285 379132
rect 550219 379067 550285 379068
rect 523794 372000 524414 378000
rect 527514 372000 528134 378000
rect 531234 372000 531854 378000
rect 534954 372000 535574 378000
rect 541794 372000 542414 378000
rect 545514 372000 546134 378000
rect 549234 372000 549854 378000
rect 520043 371924 520109 371925
rect 520043 371860 520044 371924
rect 520108 371860 520109 371924
rect 520043 371859 520109 371860
rect 549299 370972 549365 370973
rect 549299 370908 549300 370972
rect 549364 370908 549365 370972
rect 549299 370907 549365 370908
rect 518755 370836 518821 370837
rect 518755 370772 518756 370836
rect 518820 370772 518821 370836
rect 518755 370771 518821 370772
rect 518571 370564 518637 370565
rect 518571 370500 518572 370564
rect 518636 370500 518637 370564
rect 518571 370499 518637 370500
rect 454208 363454 454528 363486
rect 454208 363218 454250 363454
rect 454486 363218 454528 363454
rect 454208 363134 454528 363218
rect 454208 362898 454250 363134
rect 454486 362898 454528 363134
rect 454208 362866 454528 362898
rect 484928 363454 485248 363486
rect 484928 363218 484970 363454
rect 485206 363218 485248 363454
rect 484928 363134 485248 363218
rect 484928 362898 484970 363134
rect 485206 362898 485248 363134
rect 484928 362866 485248 362898
rect 515648 363454 515968 363486
rect 515648 363218 515690 363454
rect 515926 363218 515968 363454
rect 515648 363134 515968 363218
rect 515648 362898 515690 363134
rect 515926 362898 515968 363134
rect 515648 362866 515968 362898
rect 546368 363454 546688 363486
rect 546368 363218 546410 363454
rect 546646 363218 546688 363454
rect 546368 363134 546688 363218
rect 546368 362898 546410 363134
rect 546646 362898 546688 363134
rect 546368 362866 546688 362898
rect 469568 345454 469888 345486
rect 469568 345218 469610 345454
rect 469846 345218 469888 345454
rect 469568 345134 469888 345218
rect 469568 344898 469610 345134
rect 469846 344898 469888 345134
rect 469568 344866 469888 344898
rect 500288 345454 500608 345486
rect 500288 345218 500330 345454
rect 500566 345218 500608 345454
rect 500288 345134 500608 345218
rect 500288 344898 500330 345134
rect 500566 344898 500608 345134
rect 500288 344866 500608 344898
rect 531008 345454 531328 345486
rect 531008 345218 531050 345454
rect 531286 345218 531328 345454
rect 531008 345134 531328 345218
rect 531008 344898 531050 345134
rect 531286 344898 531328 345134
rect 531008 344866 531328 344898
rect 454208 327454 454528 327486
rect 454208 327218 454250 327454
rect 454486 327218 454528 327454
rect 454208 327134 454528 327218
rect 454208 326898 454250 327134
rect 454486 326898 454528 327134
rect 454208 326866 454528 326898
rect 484928 327454 485248 327486
rect 484928 327218 484970 327454
rect 485206 327218 485248 327454
rect 484928 327134 485248 327218
rect 484928 326898 484970 327134
rect 485206 326898 485248 327134
rect 484928 326866 485248 326898
rect 515648 327454 515968 327486
rect 515648 327218 515690 327454
rect 515926 327218 515968 327454
rect 515648 327134 515968 327218
rect 515648 326898 515690 327134
rect 515926 326898 515968 327134
rect 515648 326866 515968 326898
rect 546368 327454 546688 327486
rect 546368 327218 546410 327454
rect 546646 327218 546688 327454
rect 546368 327134 546688 327218
rect 546368 326898 546410 327134
rect 546646 326898 546688 327134
rect 546368 326866 546688 326898
rect 469568 309454 469888 309486
rect 469568 309218 469610 309454
rect 469846 309218 469888 309454
rect 469568 309134 469888 309218
rect 469568 308898 469610 309134
rect 469846 308898 469888 309134
rect 469568 308866 469888 308898
rect 500288 309454 500608 309486
rect 500288 309218 500330 309454
rect 500566 309218 500608 309454
rect 500288 309134 500608 309218
rect 500288 308898 500330 309134
rect 500566 308898 500608 309134
rect 500288 308866 500608 308898
rect 531008 309454 531328 309486
rect 531008 309218 531050 309454
rect 531286 309218 531328 309454
rect 531008 309134 531328 309218
rect 531008 308898 531050 309134
rect 531286 308898 531328 309134
rect 531008 308866 531328 308898
rect 549302 298210 549362 370907
rect 550035 370836 550101 370837
rect 550035 370772 550036 370836
rect 550100 370772 550101 370836
rect 550035 370771 550101 370772
rect 548934 298150 549362 298210
rect 451043 297804 451109 297805
rect 451043 297740 451044 297804
rect 451108 297740 451109 297804
rect 451043 297739 451109 297740
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 273454 452414 298000
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 277174 456134 298000
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 280894 459854 298000
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 284614 463574 298000
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 291454 470414 298000
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 295174 474134 298000
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 262894 477854 298000
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 266614 481574 298000
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 273454 488414 298000
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 277174 492134 298000
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 280894 495854 298000
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 284614 499574 298000
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 291454 506414 298000
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 295174 510134 298000
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 262894 513854 298000
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 266614 517574 298000
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 273454 524414 298000
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 277174 528134 298000
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 280894 531854 298000
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 284614 535574 298000
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 291454 542414 298000
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 295174 546134 298000
rect 548934 297533 548994 298150
rect 548931 297532 548997 297533
rect 548931 297468 548932 297532
rect 548996 297468 548997 297532
rect 548931 297467 548997 297468
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 262894 549854 298000
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 550038 46885 550098 370771
rect 550222 297669 550282 379067
rect 550403 378996 550469 378997
rect 550403 378932 550404 378996
rect 550468 378932 550469 378996
rect 550403 378931 550469 378932
rect 550219 297668 550285 297669
rect 550219 297604 550220 297668
rect 550284 297604 550285 297668
rect 550219 297603 550285 297604
rect 550406 297261 550466 378931
rect 550587 378860 550653 378861
rect 550587 378796 550588 378860
rect 550652 378796 550653 378860
rect 550587 378795 550653 378796
rect 550590 297805 550650 378795
rect 550771 378724 550837 378725
rect 550771 378660 550772 378724
rect 550836 378660 550837 378724
rect 550771 378659 550837 378660
rect 550774 297941 550834 378659
rect 552954 374614 553574 378000
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 550955 370700 551021 370701
rect 550955 370636 550956 370700
rect 551020 370636 551021 370700
rect 550955 370635 551021 370636
rect 550771 297940 550837 297941
rect 550771 297876 550772 297940
rect 550836 297876 550837 297940
rect 550771 297875 550837 297876
rect 550587 297804 550653 297805
rect 550587 297740 550588 297804
rect 550652 297740 550653 297804
rect 550587 297739 550653 297740
rect 550958 297397 551018 370635
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 550955 297396 551021 297397
rect 550955 297332 550956 297396
rect 551020 297332 551021 297396
rect 550955 297331 551021 297332
rect 550403 297260 550469 297261
rect 550403 297196 550404 297260
rect 550468 297196 550469 297260
rect 550403 297195 550469 297196
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 550035 46884 550101 46885
rect 550035 46820 550036 46884
rect 550100 46820 550101 46884
rect 550035 46819 550101 46820
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 558870 5677 558930 419867
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 559794 345454 560414 378000
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 558867 5676 558933 5677
rect 558867 5612 558868 5676
rect 558932 5612 558933 5676
rect 558867 5611 558933 5612
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 84250 183218 84486 183454
rect 84250 182898 84486 183134
rect 114970 183218 115206 183454
rect 114970 182898 115206 183134
rect 145690 183218 145926 183454
rect 145690 182898 145926 183134
rect 176410 183218 176646 183454
rect 176410 182898 176646 183134
rect 207130 183218 207366 183454
rect 207130 182898 207366 183134
rect 237850 183218 238086 183454
rect 237850 182898 238086 183134
rect 99610 165218 99846 165454
rect 99610 164898 99846 165134
rect 130330 165218 130566 165454
rect 130330 164898 130566 165134
rect 161050 165218 161286 165454
rect 161050 164898 161286 165134
rect 191770 165218 192006 165454
rect 191770 164898 192006 165134
rect 222490 165218 222726 165454
rect 222490 164898 222726 165134
rect 253210 165218 253446 165454
rect 253210 164898 253446 165134
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 84250 147218 84486 147454
rect 84250 146898 84486 147134
rect 114970 147218 115206 147454
rect 114970 146898 115206 147134
rect 145690 147218 145926 147454
rect 145690 146898 145926 147134
rect 176410 147218 176646 147454
rect 176410 146898 176646 147134
rect 207130 147218 207366 147454
rect 207130 146898 207366 147134
rect 237850 147218 238086 147454
rect 237850 146898 238086 147134
rect 99610 129218 99846 129454
rect 99610 128898 99846 129134
rect 130330 129218 130566 129454
rect 130330 128898 130566 129134
rect 161050 129218 161286 129454
rect 161050 128898 161286 129134
rect 191770 129218 192006 129454
rect 191770 128898 192006 129134
rect 222490 129218 222726 129454
rect 222490 128898 222726 129134
rect 253210 129218 253446 129454
rect 253210 128898 253446 129134
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 84250 111218 84486 111454
rect 84250 110898 84486 111134
rect 114970 111218 115206 111454
rect 114970 110898 115206 111134
rect 145690 111218 145926 111454
rect 145690 110898 145926 111134
rect 176410 111218 176646 111454
rect 176410 110898 176646 111134
rect 207130 111218 207366 111454
rect 207130 110898 207366 111134
rect 237850 111218 238086 111454
rect 237850 110898 238086 111134
rect 99610 93218 99846 93454
rect 99610 92898 99846 93134
rect 130330 93218 130566 93454
rect 130330 92898 130566 93134
rect 161050 93218 161286 93454
rect 161050 92898 161286 93134
rect 191770 93218 192006 93454
rect 191770 92898 192006 93134
rect 222490 93218 222726 93454
rect 222490 92898 222726 93134
rect 253210 93218 253446 93454
rect 253210 92898 253446 93134
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 539610 417218 539846 417454
rect 539610 416898 539846 417134
rect 524250 399218 524486 399454
rect 524250 398898 524486 399134
rect 554970 399218 555206 399454
rect 554970 398898 555206 399134
rect 454250 363218 454486 363454
rect 454250 362898 454486 363134
rect 484970 363218 485206 363454
rect 484970 362898 485206 363134
rect 515690 363218 515926 363454
rect 515690 362898 515926 363134
rect 546410 363218 546646 363454
rect 546410 362898 546646 363134
rect 469610 345218 469846 345454
rect 469610 344898 469846 345134
rect 500330 345218 500566 345454
rect 500330 344898 500566 345134
rect 531050 345218 531286 345454
rect 531050 344898 531286 345134
rect 454250 327218 454486 327454
rect 454250 326898 454486 327134
rect 484970 327218 485206 327454
rect 484970 326898 485206 327134
rect 515690 327218 515926 327454
rect 515690 326898 515926 327134
rect 546410 327218 546646 327454
rect 546410 326898 546646 327134
rect 469610 309218 469846 309454
rect 469610 308898 469846 309134
rect 500330 309218 500566 309454
rect 500330 308898 500566 309134
rect 531050 309218 531286 309454
rect 531050 308898 531286 309134
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 539610 417454
rect 539846 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 539610 417134
rect 539846 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 524250 399454
rect 524486 399218 554970 399454
rect 555206 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 524250 399134
rect 524486 398898 554970 399134
rect 555206 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 454250 363454
rect 454486 363218 484970 363454
rect 485206 363218 515690 363454
rect 515926 363218 546410 363454
rect 546646 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 454250 363134
rect 454486 362898 484970 363134
rect 485206 362898 515690 363134
rect 515926 362898 546410 363134
rect 546646 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 469610 345454
rect 469846 345218 500330 345454
rect 500566 345218 531050 345454
rect 531286 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 469610 345134
rect 469846 344898 500330 345134
rect 500566 344898 531050 345134
rect 531286 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 454250 327454
rect 454486 327218 484970 327454
rect 485206 327218 515690 327454
rect 515926 327218 546410 327454
rect 546646 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 454250 327134
rect 454486 326898 484970 327134
rect 485206 326898 515690 327134
rect 515926 326898 546410 327134
rect 546646 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 469610 309454
rect 469846 309218 500330 309454
rect 500566 309218 531050 309454
rect 531286 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 469610 309134
rect 469846 308898 500330 309134
rect 500566 308898 531050 309134
rect 531286 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 84250 183454
rect 84486 183218 114970 183454
rect 115206 183218 145690 183454
rect 145926 183218 176410 183454
rect 176646 183218 207130 183454
rect 207366 183218 237850 183454
rect 238086 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 84250 183134
rect 84486 182898 114970 183134
rect 115206 182898 145690 183134
rect 145926 182898 176410 183134
rect 176646 182898 207130 183134
rect 207366 182898 237850 183134
rect 238086 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 99610 165454
rect 99846 165218 130330 165454
rect 130566 165218 161050 165454
rect 161286 165218 191770 165454
rect 192006 165218 222490 165454
rect 222726 165218 253210 165454
rect 253446 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 99610 165134
rect 99846 164898 130330 165134
rect 130566 164898 161050 165134
rect 161286 164898 191770 165134
rect 192006 164898 222490 165134
rect 222726 164898 253210 165134
rect 253446 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 84250 147454
rect 84486 147218 114970 147454
rect 115206 147218 145690 147454
rect 145926 147218 176410 147454
rect 176646 147218 207130 147454
rect 207366 147218 237850 147454
rect 238086 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 84250 147134
rect 84486 146898 114970 147134
rect 115206 146898 145690 147134
rect 145926 146898 176410 147134
rect 176646 146898 207130 147134
rect 207366 146898 237850 147134
rect 238086 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 99610 129454
rect 99846 129218 130330 129454
rect 130566 129218 161050 129454
rect 161286 129218 191770 129454
rect 192006 129218 222490 129454
rect 222726 129218 253210 129454
rect 253446 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 99610 129134
rect 99846 128898 130330 129134
rect 130566 128898 161050 129134
rect 161286 128898 191770 129134
rect 192006 128898 222490 129134
rect 222726 128898 253210 129134
rect 253446 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 84250 111454
rect 84486 111218 114970 111454
rect 115206 111218 145690 111454
rect 145926 111218 176410 111454
rect 176646 111218 207130 111454
rect 207366 111218 237850 111454
rect 238086 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 84250 111134
rect 84486 110898 114970 111134
rect 115206 110898 145690 111134
rect 145926 110898 176410 111134
rect 176646 110898 207130 111134
rect 207366 110898 237850 111134
rect 238086 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 99610 93454
rect 99846 93218 130330 93454
rect 130566 93218 161050 93454
rect 161286 93218 191770 93454
rect 192006 93218 222490 93454
rect 222726 93218 253210 93454
rect 253446 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 99610 93134
rect 99846 92898 130330 93134
rect 130566 92898 161050 93134
rect 161286 92898 191770 93134
rect 192006 92898 222490 93134
rect 222726 92898 253210 93134
rect 253446 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use IOMultiplexer  ioMux
timestamp 0
transform 1 0 520000 0 1 380000
box 0 0 40000 40000
use user_proj_example  mprj
timestamp 0
transform 1 0 80000 0 1 80000
box 13 0 179846 120000
use PWM  pwm
timestamp 0
transform 1 0 450000 0 1 300000
box 0 0 100000 69080
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 78000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 78000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 78000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 78000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 78000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 372000 542414 378000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 202000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 202000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 202000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 202000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 202000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 372000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 372000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 422000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 78000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 78000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 78000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 78000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 78000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 78000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 372000 546134 378000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 202000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 202000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 202000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 202000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 202000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 202000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 372000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 372000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 422000 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 78000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 78000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 78000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 78000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 78000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 78000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 372000 549854 378000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 202000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 202000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 202000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 202000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 202000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 202000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 372000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 372000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 422000 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 78000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 78000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 78000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 78000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 78000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 378000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 202000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 202000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 202000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 202000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 202000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 372000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 372000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 422000 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 78000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 78000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 78000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 78000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 78000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 372000 531854 378000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 202000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 202000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 202000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 202000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 202000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 372000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 372000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 422000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 78000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 78000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 78000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 78000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 78000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 372000 535574 378000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 202000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 202000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 202000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 202000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 202000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 372000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 372000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 422000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 78000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 78000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 78000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 78000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 78000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 372000 524414 378000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 378000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 202000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 202000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 202000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 202000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 202000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 372000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 372000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 422000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 422000 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 78000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 78000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 78000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 78000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 78000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 372000 528134 378000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 202000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 202000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 202000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 202000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 202000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 372000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 372000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 422000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
