VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Art
  CLASS BLOCK ;
  FOREIGN Art ;
  ORIGIN -0.200 0.000 ;
  SIZE 753.320 BY 300.000 ;
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.20000 0.00000 1.00000 300.00000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 749.00000 0.00000 749.80000 300.00000 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.000 30.000 105.000 70.000 ;
        RECT 5.000 5.000 25.000 25.000 ;
      LAYER met1 ;
        RECT 85.000 60.000 105.000 70.120 ;
        RECT 65.000 50.000 105.000 60.000 ;
        RECT 45.000 40.000 105.000 50.000 ;
        RECT 25.000 30.120 105.000 40.000 ;
        RECT 25.000 30.000 85.000 30.120 ;
        RECT 25.000 5.000 45.000 25.000 ;
      LAYER met2 ;
        RECT 45.000 60.000 65.000 70.000 ;
        RECT 25.000 50.000 45.000 60.000 ;
        RECT 85.000 50.000 105.000 60.000 ;
        RECT 5.000 40.000 25.000 50.000 ;
        RECT 65.000 40.000 105.000 50.000 ;
        RECT 45.000 30.000 105.000 40.000 ;
        RECT 45.000 5.000 65.000 25.000 ;
      LAYER met3 ;
        RECT 25.000 60.000 45.000 70.000 ;
        RECT 5.000 50.000 25.000 60.000 ;
        RECT 85.000 40.000 105.000 50.000 ;
        RECT 65.000 30.000 105.000 40.000 ;
        RECT 65.000 5.000 85.000 25.000 ;
      LAYER met4 ;
        RECT 0.200 0.000 1.000 300.000 ;
        RECT 369.830 289.290 375.830 291.290 ;
        RECT 369.830 287.290 371.830 289.290 ;
        RECT 367.830 285.290 371.830 287.290 ;
        RECT 373.830 287.290 375.830 289.290 ;
        RECT 519.830 289.290 525.830 291.290 ;
        RECT 519.830 287.290 521.830 289.290 ;
        RECT 373.830 285.290 377.830 287.290 ;
        RECT 367.830 281.290 369.830 285.290 ;
        RECT 365.830 279.290 369.830 281.290 ;
        RECT 375.830 281.290 377.830 285.290 ;
        RECT 517.830 285.290 521.830 287.290 ;
        RECT 523.830 287.290 525.830 289.290 ;
        RECT 669.830 289.290 675.830 291.290 ;
        RECT 669.830 287.290 671.830 289.290 ;
        RECT 523.830 285.290 527.830 287.290 ;
        RECT 517.830 281.290 519.830 285.290 ;
        RECT 375.830 279.290 379.830 281.290 ;
        RECT 365.830 275.290 367.830 279.290 ;
        RECT 363.830 273.290 367.830 275.290 ;
        RECT 369.830 273.290 373.830 277.290 ;
        RECT 377.830 275.290 379.830 279.290 ;
        RECT 515.830 279.290 519.830 281.290 ;
        RECT 525.830 281.290 527.830 285.290 ;
        RECT 667.830 285.290 671.830 287.290 ;
        RECT 673.830 287.290 675.830 289.290 ;
        RECT 673.830 285.290 677.830 287.290 ;
        RECT 667.830 281.290 669.830 285.290 ;
        RECT 525.830 279.290 529.830 281.290 ;
        RECT 515.830 275.290 517.830 279.290 ;
        RECT 377.830 273.290 381.830 275.290 ;
        RECT 363.830 269.290 365.830 273.290 ;
        RECT 361.830 267.290 365.830 269.290 ;
        RECT 367.830 271.290 373.830 273.290 ;
        RECT 379.830 271.290 381.830 273.290 ;
        RECT 513.830 273.290 517.830 275.290 ;
        RECT 519.830 273.290 523.830 277.290 ;
        RECT 527.830 275.290 529.830 279.290 ;
        RECT 665.830 279.290 669.830 281.290 ;
        RECT 675.830 281.290 677.830 285.290 ;
        RECT 675.830 279.290 679.830 281.290 ;
        RECT 665.830 275.290 667.830 279.290 ;
        RECT 527.830 273.290 531.830 275.290 ;
        RECT 367.830 269.290 375.830 271.290 ;
        RECT 379.830 269.290 383.830 271.290 ;
        RECT 513.830 269.290 515.830 273.290 ;
        RECT 367.830 267.290 377.830 269.290 ;
        RECT 361.830 265.290 363.830 267.290 ;
        RECT 359.830 263.290 363.830 265.290 ;
        RECT 365.830 263.290 373.830 267.290 ;
        RECT 359.830 259.290 361.830 263.290 ;
        RECT 357.830 257.290 361.830 259.290 ;
        RECT 363.830 259.290 373.830 263.290 ;
        RECT 375.830 263.290 379.830 267.290 ;
        RECT 381.830 265.290 383.830 269.290 ;
        RECT 511.830 267.290 515.830 269.290 ;
        RECT 517.830 271.290 523.830 273.290 ;
        RECT 529.830 271.290 531.830 273.290 ;
        RECT 663.830 273.290 667.830 275.290 ;
        RECT 669.830 273.290 673.830 277.290 ;
        RECT 677.830 275.290 679.830 279.290 ;
        RECT 677.830 273.290 681.830 275.290 ;
        RECT 517.830 269.290 525.830 271.290 ;
        RECT 529.830 269.290 533.830 271.290 ;
        RECT 663.830 269.290 665.830 273.290 ;
        RECT 517.830 267.290 527.830 269.290 ;
        RECT 511.830 265.290 513.830 267.290 ;
        RECT 381.830 263.290 385.830 265.290 ;
        RECT 375.830 259.290 381.830 263.290 ;
        RECT 363.830 257.290 375.830 259.290 ;
        RECT 357.830 255.290 359.830 257.290 ;
        RECT 351.830 253.290 359.830 255.290 ;
        RECT 361.830 253.290 375.830 257.290 ;
        RECT 377.830 257.290 381.830 259.290 ;
        RECT 383.830 259.290 385.830 263.290 ;
        RECT 509.830 263.290 513.830 265.290 ;
        RECT 515.830 263.290 523.830 267.290 ;
        RECT 509.830 259.290 511.830 263.290 ;
        RECT 383.830 257.290 387.830 259.290 ;
        RECT 377.830 255.290 383.830 257.290 ;
        RECT 377.830 253.290 379.830 255.290 ;
        RECT 385.830 253.290 387.830 257.290 ;
        RECT 507.830 257.290 511.830 259.290 ;
        RECT 513.830 259.290 523.830 263.290 ;
        RECT 525.830 263.290 529.830 267.290 ;
        RECT 531.830 265.290 533.830 269.290 ;
        RECT 661.830 267.290 665.830 269.290 ;
        RECT 667.830 271.290 673.830 273.290 ;
        RECT 679.830 271.290 681.830 273.290 ;
        RECT 667.830 269.290 675.830 271.290 ;
        RECT 679.830 269.290 683.830 271.290 ;
        RECT 667.830 267.290 677.830 269.290 ;
        RECT 661.830 265.290 663.830 267.290 ;
        RECT 531.830 263.290 535.830 265.290 ;
        RECT 525.830 259.290 531.830 263.290 ;
        RECT 513.830 257.290 525.830 259.290 ;
        RECT 507.830 255.290 509.830 257.290 ;
        RECT 501.830 253.290 509.830 255.290 ;
        RECT 511.830 253.290 525.830 257.290 ;
        RECT 527.830 257.290 531.830 259.290 ;
        RECT 533.830 259.290 535.830 263.290 ;
        RECT 659.830 263.290 663.830 265.290 ;
        RECT 665.830 263.290 673.830 267.290 ;
        RECT 659.830 259.290 661.830 263.290 ;
        RECT 533.830 257.290 537.830 259.290 ;
        RECT 527.830 255.290 533.830 257.290 ;
        RECT 527.830 253.290 529.830 255.290 ;
        RECT 535.830 253.290 537.830 257.290 ;
        RECT 657.830 257.290 661.830 259.290 ;
        RECT 663.830 259.290 673.830 263.290 ;
        RECT 675.830 263.290 679.830 267.290 ;
        RECT 681.830 265.290 683.830 269.290 ;
        RECT 681.830 263.290 685.830 265.290 ;
        RECT 675.830 259.290 681.830 263.290 ;
        RECT 663.830 257.290 675.830 259.290 ;
        RECT 657.830 255.290 659.830 257.290 ;
        RECT 651.830 253.290 659.830 255.290 ;
        RECT 661.830 253.290 675.830 257.290 ;
        RECT 677.830 257.290 681.830 259.290 ;
        RECT 683.830 259.290 685.830 263.290 ;
        RECT 683.830 257.290 687.830 259.290 ;
        RECT 677.830 255.290 683.830 257.290 ;
        RECT 677.830 253.290 679.830 255.290 ;
        RECT 685.830 253.290 687.830 257.290 ;
        RECT 341.830 251.290 353.830 253.290 ;
        RECT 361.830 251.290 377.830 253.290 ;
        RECT 379.830 251.290 383.830 253.290 ;
        RECT 385.830 251.290 395.830 253.290 ;
        RECT 491.830 251.290 503.830 253.290 ;
        RECT 511.830 251.290 527.830 253.290 ;
        RECT 529.830 251.290 533.830 253.290 ;
        RECT 535.830 251.290 545.830 253.290 ;
        RECT 641.830 251.290 653.830 253.290 ;
        RECT 661.830 251.290 677.830 253.290 ;
        RECT 679.830 251.290 683.830 253.290 ;
        RECT 685.830 251.290 695.830 253.290 ;
        RECT 335.830 249.290 343.830 251.290 ;
        RECT 353.830 249.290 357.830 251.290 ;
        RECT 335.830 245.290 337.830 249.290 ;
        RECT 343.830 247.290 357.830 249.290 ;
        RECT 359.830 247.290 385.830 251.290 ;
        RECT 393.830 249.290 403.830 251.290 ;
        RECT 485.830 249.290 493.830 251.290 ;
        RECT 503.830 249.290 507.830 251.290 ;
        RECT 387.830 247.290 389.830 249.290 ;
        RECT 401.830 247.290 411.830 249.290 ;
        RECT 343.830 245.290 359.830 247.290 ;
        RECT 369.830 245.290 381.830 247.290 ;
        RECT 385.830 245.290 393.830 247.290 ;
        RECT 409.830 245.290 415.830 247.290 ;
        RECT 335.830 243.290 343.830 245.290 ;
        RECT 353.830 243.290 369.830 245.290 ;
        RECT 381.830 243.290 399.830 245.290 ;
        RECT 413.830 243.290 415.830 245.290 ;
        RECT 485.830 245.290 487.830 249.290 ;
        RECT 493.830 247.290 507.830 249.290 ;
        RECT 509.830 247.290 535.830 251.290 ;
        RECT 543.830 249.290 553.830 251.290 ;
        RECT 635.830 249.290 643.830 251.290 ;
        RECT 653.830 249.290 657.830 251.290 ;
        RECT 537.830 247.290 539.830 249.290 ;
        RECT 551.830 247.290 561.830 249.290 ;
        RECT 493.830 245.290 509.830 247.290 ;
        RECT 519.830 245.290 531.830 247.290 ;
        RECT 535.830 245.290 543.830 247.290 ;
        RECT 559.830 245.290 565.830 247.290 ;
        RECT 485.830 243.290 493.830 245.290 ;
        RECT 503.830 243.290 519.830 245.290 ;
        RECT 531.830 243.290 549.830 245.290 ;
        RECT 563.830 243.290 565.830 245.290 ;
        RECT 635.830 245.290 637.830 249.290 ;
        RECT 643.830 247.290 657.830 249.290 ;
        RECT 659.830 247.290 685.830 251.290 ;
        RECT 693.830 249.290 703.830 251.290 ;
        RECT 687.830 247.290 689.830 249.290 ;
        RECT 701.830 247.290 711.830 249.290 ;
        RECT 643.830 245.290 659.830 247.290 ;
        RECT 669.830 245.290 681.830 247.290 ;
        RECT 685.830 245.290 693.830 247.290 ;
        RECT 709.830 245.290 715.830 247.290 ;
        RECT 635.830 243.290 643.830 245.290 ;
        RECT 653.830 243.290 669.830 245.290 ;
        RECT 681.830 243.290 699.830 245.290 ;
        RECT 713.830 243.290 715.830 245.290 ;
        RECT 341.830 241.290 353.830 243.290 ;
        RECT 363.830 241.290 403.830 243.290 ;
        RECT 411.830 241.290 415.830 243.290 ;
        RECT 491.830 241.290 503.830 243.290 ;
        RECT 513.830 241.290 553.830 243.290 ;
        RECT 561.830 241.290 565.830 243.290 ;
        RECT 641.830 241.290 653.830 243.290 ;
        RECT 663.830 241.290 703.830 243.290 ;
        RECT 711.830 241.290 715.830 243.290 ;
        RECT 351.830 239.290 363.830 241.290 ;
        RECT 373.830 239.290 401.830 241.290 ;
        RECT 409.830 239.290 413.830 241.290 ;
        RECT 501.830 239.290 513.830 241.290 ;
        RECT 523.830 239.290 551.830 241.290 ;
        RECT 559.830 239.290 563.830 241.290 ;
        RECT 651.830 239.290 663.830 241.290 ;
        RECT 673.830 239.290 701.830 241.290 ;
        RECT 709.830 239.290 713.830 241.290 ;
        RECT 353.830 237.290 355.830 239.290 ;
        RECT 351.830 235.290 355.830 237.290 ;
        RECT 357.830 237.290 373.830 239.290 ;
        RECT 383.830 237.290 393.830 239.290 ;
        RECT 401.830 237.290 411.830 239.290 ;
        RECT 503.830 237.290 505.830 239.290 ;
        RECT 357.830 235.290 383.830 237.290 ;
        RECT 393.830 235.290 403.830 237.290 ;
        RECT 501.830 235.290 505.830 237.290 ;
        RECT 507.830 237.290 523.830 239.290 ;
        RECT 533.830 237.290 543.830 239.290 ;
        RECT 551.830 237.290 561.830 239.290 ;
        RECT 653.830 237.290 655.830 239.290 ;
        RECT 507.830 235.290 533.830 237.290 ;
        RECT 543.830 235.290 553.830 237.290 ;
        RECT 651.830 235.290 655.830 237.290 ;
        RECT 657.830 237.290 673.830 239.290 ;
        RECT 683.830 237.290 693.830 239.290 ;
        RECT 701.830 237.290 711.830 239.290 ;
        RECT 657.830 235.290 683.830 237.290 ;
        RECT 693.830 235.290 703.830 237.290 ;
        RECT 351.830 229.290 353.830 235.290 ;
        RECT 355.830 233.290 373.830 235.290 ;
        RECT 383.830 233.290 395.830 235.290 ;
        RECT 355.830 231.290 371.830 233.290 ;
        RECT 357.830 229.290 371.830 231.290 ;
        RECT 373.830 231.290 377.830 233.290 ;
        RECT 381.830 231.290 383.830 233.290 ;
        RECT 387.830 231.290 389.830 233.290 ;
        RECT 393.830 231.290 395.830 233.290 ;
        RECT 403.830 231.290 409.830 233.290 ;
        RECT 373.830 229.290 375.830 231.290 ;
        RECT 387.830 229.290 395.830 231.290 ;
        RECT 401.830 229.290 405.830 231.290 ;
        RECT 407.830 229.290 409.830 231.290 ;
        RECT 501.830 229.290 503.830 235.290 ;
        RECT 505.830 233.290 523.830 235.290 ;
        RECT 533.830 233.290 545.830 235.290 ;
        RECT 505.830 231.290 521.830 233.290 ;
        RECT 507.830 229.290 521.830 231.290 ;
        RECT 523.830 231.290 527.830 233.290 ;
        RECT 531.830 231.290 533.830 233.290 ;
        RECT 537.830 231.290 539.830 233.290 ;
        RECT 543.830 231.290 545.830 233.290 ;
        RECT 553.830 231.290 559.830 233.290 ;
        RECT 523.830 229.290 525.830 231.290 ;
        RECT 537.830 229.290 545.830 231.290 ;
        RECT 551.830 229.290 555.830 231.290 ;
        RECT 557.830 229.290 559.830 231.290 ;
        RECT 651.830 229.290 653.830 235.290 ;
        RECT 655.830 233.290 673.830 235.290 ;
        RECT 683.830 233.290 695.830 235.290 ;
        RECT 655.830 231.290 671.830 233.290 ;
        RECT 657.830 229.290 671.830 231.290 ;
        RECT 673.830 231.290 677.830 233.290 ;
        RECT 681.830 231.290 683.830 233.290 ;
        RECT 687.830 231.290 689.830 233.290 ;
        RECT 693.830 231.290 695.830 233.290 ;
        RECT 703.830 231.290 709.830 233.290 ;
        RECT 673.830 229.290 675.830 231.290 ;
        RECT 687.830 229.290 695.830 231.290 ;
        RECT 701.830 229.290 705.830 231.290 ;
        RECT 707.830 229.290 709.830 231.290 ;
        RECT 349.830 227.290 355.830 229.290 ;
        RECT 347.830 225.290 351.830 227.290 ;
        RECT 353.830 225.290 359.830 227.290 ;
        RECT 361.830 225.290 371.830 229.290 ;
        RECT 375.830 227.290 377.830 229.290 ;
        RECT 387.830 227.290 391.830 229.290 ;
        RECT 397.830 227.290 403.830 229.290 ;
        RECT 405.830 227.290 409.830 229.290 ;
        RECT 499.830 227.290 505.830 229.290 ;
        RECT 385.830 225.290 391.830 227.290 ;
        RECT 393.830 225.290 399.830 227.290 ;
        RECT 345.830 223.290 349.830 225.290 ;
        RECT 351.830 223.290 361.830 225.290 ;
        RECT 365.830 223.290 373.830 225.290 ;
        RECT 379.830 223.290 395.830 225.290 ;
        RECT 399.830 223.290 403.830 225.290 ;
        RECT 345.830 217.290 347.830 223.290 ;
        RECT 343.830 215.290 347.830 217.290 ;
        RECT 349.830 221.290 363.830 223.290 ;
        RECT 367.830 221.290 373.830 223.290 ;
        RECT 383.830 221.290 391.830 223.290 ;
        RECT 395.830 221.290 405.830 223.290 ;
        RECT 407.830 221.290 409.830 227.290 ;
        RECT 497.830 225.290 501.830 227.290 ;
        RECT 503.830 225.290 509.830 227.290 ;
        RECT 511.830 225.290 521.830 229.290 ;
        RECT 525.830 227.290 527.830 229.290 ;
        RECT 537.830 227.290 541.830 229.290 ;
        RECT 547.830 227.290 553.830 229.290 ;
        RECT 555.830 227.290 559.830 229.290 ;
        RECT 649.830 227.290 655.830 229.290 ;
        RECT 535.830 225.290 541.830 227.290 ;
        RECT 543.830 225.290 549.830 227.290 ;
        RECT 349.830 219.290 367.830 221.290 ;
        RECT 369.830 219.290 373.830 221.290 ;
        RECT 381.830 219.290 387.830 221.290 ;
        RECT 391.830 219.290 401.830 221.290 ;
        RECT 405.830 219.290 409.830 221.290 ;
        RECT 495.830 223.290 499.830 225.290 ;
        RECT 501.830 223.290 511.830 225.290 ;
        RECT 515.830 223.290 523.830 225.290 ;
        RECT 529.830 223.290 545.830 225.290 ;
        RECT 549.830 223.290 553.830 225.290 ;
        RECT 349.830 217.290 369.830 219.290 ;
        RECT 377.830 217.290 383.830 219.290 ;
        RECT 387.830 217.290 399.830 219.290 ;
        RECT 349.830 215.290 389.830 217.290 ;
        RECT 397.830 215.290 399.830 217.290 ;
        RECT 401.830 217.290 407.830 219.290 ;
        RECT 495.830 217.290 497.830 223.290 ;
        RECT 401.830 215.290 403.830 217.290 ;
        RECT 343.830 195.290 345.830 215.290 ;
        RECT 347.830 213.290 363.830 215.290 ;
        RECT 365.830 213.290 367.830 215.290 ;
        RECT 371.830 213.290 383.830 215.290 ;
        RECT 347.830 211.290 361.830 213.290 ;
        RECT 363.830 211.290 365.830 213.290 ;
        RECT 367.830 211.290 371.830 213.290 ;
        RECT 377.830 211.290 381.830 213.290 ;
        RECT 383.830 211.290 385.830 213.290 ;
        RECT 399.830 211.290 403.830 215.290 ;
        RECT 347.830 209.290 363.830 211.290 ;
        RECT 365.830 209.290 367.830 211.290 ;
        RECT 347.830 207.290 361.830 209.290 ;
        RECT 363.830 207.290 367.830 209.290 ;
        RECT 371.830 209.290 381.830 211.290 ;
        RECT 385.830 209.290 403.830 211.290 ;
        RECT 493.830 215.290 497.830 217.290 ;
        RECT 499.830 221.290 513.830 223.290 ;
        RECT 517.830 221.290 523.830 223.290 ;
        RECT 533.830 221.290 541.830 223.290 ;
        RECT 545.830 221.290 555.830 223.290 ;
        RECT 557.830 221.290 559.830 227.290 ;
        RECT 647.830 225.290 651.830 227.290 ;
        RECT 653.830 225.290 659.830 227.290 ;
        RECT 661.830 225.290 671.830 229.290 ;
        RECT 675.830 227.290 677.830 229.290 ;
        RECT 687.830 227.290 691.830 229.290 ;
        RECT 697.830 227.290 703.830 229.290 ;
        RECT 705.830 227.290 709.830 229.290 ;
        RECT 685.830 225.290 691.830 227.290 ;
        RECT 693.830 225.290 699.830 227.290 ;
        RECT 499.830 219.290 517.830 221.290 ;
        RECT 519.830 219.290 523.830 221.290 ;
        RECT 531.830 219.290 537.830 221.290 ;
        RECT 541.830 219.290 551.830 221.290 ;
        RECT 555.830 219.290 559.830 221.290 ;
        RECT 645.830 223.290 649.830 225.290 ;
        RECT 651.830 223.290 661.830 225.290 ;
        RECT 665.830 223.290 673.830 225.290 ;
        RECT 679.830 223.290 695.830 225.290 ;
        RECT 699.830 223.290 703.830 225.290 ;
        RECT 499.830 217.290 519.830 219.290 ;
        RECT 527.830 217.290 533.830 219.290 ;
        RECT 537.830 217.290 549.830 219.290 ;
        RECT 499.830 215.290 539.830 217.290 ;
        RECT 547.830 215.290 549.830 217.290 ;
        RECT 551.830 217.290 557.830 219.290 ;
        RECT 645.830 217.290 647.830 223.290 ;
        RECT 551.830 215.290 553.830 217.290 ;
        RECT 371.830 207.290 373.830 209.290 ;
        RECT 379.830 207.290 383.830 209.290 ;
        RECT 387.830 207.290 389.830 209.290 ;
        RECT 401.830 207.290 405.830 209.290 ;
        RECT 347.830 205.290 363.830 207.290 ;
        RECT 365.830 205.290 367.830 207.290 ;
        RECT 373.830 205.290 377.830 207.290 ;
        RECT 347.830 203.290 365.830 205.290 ;
        RECT 367.830 203.290 369.830 205.290 ;
        RECT 375.830 203.290 377.830 205.290 ;
        RECT 379.830 205.290 381.830 207.290 ;
        RECT 379.830 203.290 383.830 205.290 ;
        RECT 385.830 203.290 387.830 207.290 ;
        RECT 403.830 205.290 407.830 207.290 ;
        RECT 399.830 203.290 403.830 205.290 ;
        RECT 347.830 201.290 363.830 203.290 ;
        RECT 369.830 201.290 371.830 203.290 ;
        RECT 377.830 201.290 385.830 203.290 ;
        RECT 387.830 201.290 391.830 203.290 ;
        RECT 395.830 201.290 401.830 203.290 ;
        RECT 405.830 201.290 407.830 205.290 ;
        RECT 347.830 199.290 365.830 201.290 ;
        RECT 371.830 199.290 373.830 201.290 ;
        RECT 381.830 199.290 387.830 201.290 ;
        RECT 391.830 199.290 395.830 201.290 ;
        RECT 401.830 199.290 407.830 201.290 ;
        RECT 347.830 197.290 363.830 199.290 ;
        RECT 373.830 197.290 375.830 199.290 ;
        RECT 383.830 197.290 391.830 199.290 ;
        RECT 395.830 197.290 403.830 199.290 ;
        RECT 347.830 195.290 361.830 197.290 ;
        RECT 363.830 195.290 365.830 197.290 ;
        RECT 375.830 195.290 379.830 197.290 ;
        RECT 389.830 195.290 397.830 197.290 ;
        RECT 493.830 195.290 495.830 215.290 ;
        RECT 497.830 213.290 513.830 215.290 ;
        RECT 515.830 213.290 517.830 215.290 ;
        RECT 521.830 213.290 533.830 215.290 ;
        RECT 497.830 211.290 511.830 213.290 ;
        RECT 513.830 211.290 515.830 213.290 ;
        RECT 517.830 211.290 521.830 213.290 ;
        RECT 527.830 211.290 531.830 213.290 ;
        RECT 533.830 211.290 535.830 213.290 ;
        RECT 549.830 211.290 553.830 215.290 ;
        RECT 497.830 209.290 513.830 211.290 ;
        RECT 515.830 209.290 517.830 211.290 ;
        RECT 497.830 207.290 511.830 209.290 ;
        RECT 513.830 207.290 517.830 209.290 ;
        RECT 521.830 209.290 531.830 211.290 ;
        RECT 535.830 209.290 553.830 211.290 ;
        RECT 643.830 215.290 647.830 217.290 ;
        RECT 649.830 221.290 663.830 223.290 ;
        RECT 667.830 221.290 673.830 223.290 ;
        RECT 683.830 221.290 691.830 223.290 ;
        RECT 695.830 221.290 705.830 223.290 ;
        RECT 707.830 221.290 709.830 227.290 ;
        RECT 649.830 219.290 667.830 221.290 ;
        RECT 669.830 219.290 673.830 221.290 ;
        RECT 681.830 219.290 687.830 221.290 ;
        RECT 691.830 219.290 701.830 221.290 ;
        RECT 705.830 219.290 709.830 221.290 ;
        RECT 649.830 217.290 669.830 219.290 ;
        RECT 677.830 217.290 683.830 219.290 ;
        RECT 687.830 217.290 699.830 219.290 ;
        RECT 649.830 215.290 689.830 217.290 ;
        RECT 697.830 215.290 699.830 217.290 ;
        RECT 701.830 217.290 707.830 219.290 ;
        RECT 701.830 215.290 703.830 217.290 ;
        RECT 521.830 207.290 523.830 209.290 ;
        RECT 529.830 207.290 533.830 209.290 ;
        RECT 537.830 207.290 539.830 209.290 ;
        RECT 551.830 207.290 555.830 209.290 ;
        RECT 497.830 205.290 513.830 207.290 ;
        RECT 515.830 205.290 517.830 207.290 ;
        RECT 523.830 205.290 527.830 207.290 ;
        RECT 497.830 203.290 515.830 205.290 ;
        RECT 517.830 203.290 519.830 205.290 ;
        RECT 525.830 203.290 527.830 205.290 ;
        RECT 529.830 205.290 531.830 207.290 ;
        RECT 529.830 203.290 533.830 205.290 ;
        RECT 535.830 203.290 537.830 207.290 ;
        RECT 553.830 205.290 557.830 207.290 ;
        RECT 549.830 203.290 553.830 205.290 ;
        RECT 497.830 201.290 513.830 203.290 ;
        RECT 519.830 201.290 521.830 203.290 ;
        RECT 527.830 201.290 535.830 203.290 ;
        RECT 537.830 201.290 541.830 203.290 ;
        RECT 545.830 201.290 551.830 203.290 ;
        RECT 555.830 201.290 557.830 205.290 ;
        RECT 497.830 199.290 515.830 201.290 ;
        RECT 521.830 199.290 523.830 201.290 ;
        RECT 531.830 199.290 537.830 201.290 ;
        RECT 541.830 199.290 545.830 201.290 ;
        RECT 551.830 199.290 557.830 201.290 ;
        RECT 497.830 197.290 513.830 199.290 ;
        RECT 523.830 197.290 525.830 199.290 ;
        RECT 533.830 197.290 541.830 199.290 ;
        RECT 545.830 197.290 553.830 199.290 ;
        RECT 497.830 195.290 511.830 197.290 ;
        RECT 513.830 195.290 515.830 197.290 ;
        RECT 525.830 195.290 529.830 197.290 ;
        RECT 539.830 195.290 547.830 197.290 ;
        RECT 643.830 195.290 645.830 215.290 ;
        RECT 647.830 213.290 663.830 215.290 ;
        RECT 665.830 213.290 667.830 215.290 ;
        RECT 671.830 213.290 683.830 215.290 ;
        RECT 647.830 211.290 661.830 213.290 ;
        RECT 663.830 211.290 665.830 213.290 ;
        RECT 667.830 211.290 671.830 213.290 ;
        RECT 677.830 211.290 681.830 213.290 ;
        RECT 683.830 211.290 685.830 213.290 ;
        RECT 699.830 211.290 703.830 215.290 ;
        RECT 647.830 209.290 663.830 211.290 ;
        RECT 665.830 209.290 667.830 211.290 ;
        RECT 647.830 207.290 661.830 209.290 ;
        RECT 663.830 207.290 667.830 209.290 ;
        RECT 671.830 209.290 681.830 211.290 ;
        RECT 685.830 209.290 703.830 211.290 ;
        RECT 671.830 207.290 673.830 209.290 ;
        RECT 679.830 207.290 683.830 209.290 ;
        RECT 687.830 207.290 689.830 209.290 ;
        RECT 701.830 207.290 705.830 209.290 ;
        RECT 647.830 205.290 663.830 207.290 ;
        RECT 665.830 205.290 667.830 207.290 ;
        RECT 673.830 205.290 677.830 207.290 ;
        RECT 647.830 203.290 665.830 205.290 ;
        RECT 667.830 203.290 669.830 205.290 ;
        RECT 675.830 203.290 677.830 205.290 ;
        RECT 679.830 205.290 681.830 207.290 ;
        RECT 679.830 203.290 683.830 205.290 ;
        RECT 685.830 203.290 687.830 207.290 ;
        RECT 703.830 205.290 707.830 207.290 ;
        RECT 699.830 203.290 703.830 205.290 ;
        RECT 647.830 201.290 663.830 203.290 ;
        RECT 669.830 201.290 671.830 203.290 ;
        RECT 677.830 201.290 685.830 203.290 ;
        RECT 687.830 201.290 691.830 203.290 ;
        RECT 695.830 201.290 701.830 203.290 ;
        RECT 705.830 201.290 707.830 205.290 ;
        RECT 647.830 199.290 665.830 201.290 ;
        RECT 671.830 199.290 673.830 201.290 ;
        RECT 681.830 199.290 687.830 201.290 ;
        RECT 691.830 199.290 695.830 201.290 ;
        RECT 701.830 199.290 707.830 201.290 ;
        RECT 647.830 197.290 663.830 199.290 ;
        RECT 673.830 197.290 675.830 199.290 ;
        RECT 683.830 197.290 691.830 199.290 ;
        RECT 695.830 197.290 703.830 199.290 ;
        RECT 647.830 195.290 661.830 197.290 ;
        RECT 663.830 195.290 665.830 197.290 ;
        RECT 675.830 195.290 679.830 197.290 ;
        RECT 689.830 195.290 697.830 197.290 ;
        RECT 343.830 193.290 347.830 195.290 ;
        RECT 345.830 177.290 347.830 193.290 ;
        RECT 349.830 191.290 359.830 195.290 ;
        RECT 361.830 193.290 363.830 195.290 ;
        RECT 365.830 193.290 367.830 195.290 ;
        RECT 379.830 193.290 393.830 195.290 ;
        RECT 493.830 193.290 497.830 195.290 ;
        RECT 363.830 191.290 365.830 193.290 ;
        RECT 379.830 191.290 389.830 193.290 ;
        RECT 349.830 189.290 363.830 191.290 ;
        RECT 365.830 189.290 367.830 191.290 ;
        RECT 381.830 189.290 389.830 191.290 ;
        RECT 349.830 187.290 361.830 189.290 ;
        RECT 363.830 187.290 365.830 189.290 ;
        RECT 349.830 185.290 363.830 187.290 ;
        RECT 365.830 185.290 367.830 187.290 ;
        RECT 381.830 185.290 391.830 189.290 ;
        RECT 349.830 183.290 365.830 185.290 ;
        RECT 349.830 181.290 363.830 183.290 ;
        RECT 365.830 181.290 367.830 183.290 ;
        RECT 383.830 181.290 391.830 185.290 ;
        RECT 349.830 179.290 365.830 181.290 ;
        RECT 349.830 177.290 363.830 179.290 ;
        RECT 365.830 177.290 367.830 179.290 ;
        RECT 385.830 177.290 391.830 181.290 ;
        RECT 345.830 175.290 349.830 177.290 ;
        RECT 351.830 175.290 365.830 177.290 ;
        RECT 383.830 175.290 385.830 177.290 ;
        RECT 389.830 175.290 391.830 177.290 ;
        RECT 495.830 177.290 497.830 193.290 ;
        RECT 499.830 191.290 509.830 195.290 ;
        RECT 511.830 193.290 513.830 195.290 ;
        RECT 515.830 193.290 517.830 195.290 ;
        RECT 529.830 193.290 543.830 195.290 ;
        RECT 643.830 193.290 647.830 195.290 ;
        RECT 513.830 191.290 515.830 193.290 ;
        RECT 529.830 191.290 539.830 193.290 ;
        RECT 499.830 189.290 513.830 191.290 ;
        RECT 515.830 189.290 517.830 191.290 ;
        RECT 531.830 189.290 539.830 191.290 ;
        RECT 499.830 187.290 511.830 189.290 ;
        RECT 513.830 187.290 515.830 189.290 ;
        RECT 499.830 185.290 513.830 187.290 ;
        RECT 515.830 185.290 517.830 187.290 ;
        RECT 531.830 185.290 541.830 189.290 ;
        RECT 499.830 183.290 515.830 185.290 ;
        RECT 499.830 181.290 513.830 183.290 ;
        RECT 515.830 181.290 517.830 183.290 ;
        RECT 533.830 181.290 541.830 185.290 ;
        RECT 499.830 179.290 515.830 181.290 ;
        RECT 499.830 177.290 513.830 179.290 ;
        RECT 515.830 177.290 517.830 179.290 ;
        RECT 535.830 177.290 541.830 181.290 ;
        RECT 495.830 175.290 499.830 177.290 ;
        RECT 501.830 175.290 515.830 177.290 ;
        RECT 533.830 175.290 535.830 177.290 ;
        RECT 539.830 175.290 541.830 177.290 ;
        RECT 645.830 177.290 647.830 193.290 ;
        RECT 649.830 191.290 659.830 195.290 ;
        RECT 661.830 193.290 663.830 195.290 ;
        RECT 665.830 193.290 667.830 195.290 ;
        RECT 679.830 193.290 693.830 195.290 ;
        RECT 663.830 191.290 665.830 193.290 ;
        RECT 679.830 191.290 689.830 193.290 ;
        RECT 649.830 189.290 663.830 191.290 ;
        RECT 665.830 189.290 667.830 191.290 ;
        RECT 681.830 189.290 689.830 191.290 ;
        RECT 649.830 187.290 661.830 189.290 ;
        RECT 663.830 187.290 665.830 189.290 ;
        RECT 649.830 185.290 663.830 187.290 ;
        RECT 665.830 185.290 667.830 187.290 ;
        RECT 681.830 185.290 691.830 189.290 ;
        RECT 649.830 183.290 665.830 185.290 ;
        RECT 649.830 181.290 663.830 183.290 ;
        RECT 665.830 181.290 667.830 183.290 ;
        RECT 683.830 181.290 691.830 185.290 ;
        RECT 649.830 179.290 665.830 181.290 ;
        RECT 649.830 177.290 663.830 179.290 ;
        RECT 665.830 177.290 667.830 179.290 ;
        RECT 685.830 177.290 691.830 181.290 ;
        RECT 645.830 175.290 649.830 177.290 ;
        RECT 651.830 175.290 665.830 177.290 ;
        RECT 683.830 175.290 685.830 177.290 ;
        RECT 689.830 175.290 691.830 177.290 ;
        RECT 347.830 173.290 349.830 175.290 ;
        RECT 355.830 173.290 363.830 175.290 ;
        RECT 365.830 173.290 367.830 175.290 ;
        RECT 369.830 173.290 371.830 175.290 ;
        RECT 373.830 173.290 375.830 175.290 ;
        RECT 377.830 173.290 379.830 175.290 ;
        RECT 381.830 173.290 383.830 175.290 ;
        RECT 385.830 173.290 391.830 175.290 ;
        RECT 497.830 173.290 499.830 175.290 ;
        RECT 505.830 173.290 513.830 175.290 ;
        RECT 515.830 173.290 517.830 175.290 ;
        RECT 519.830 173.290 521.830 175.290 ;
        RECT 523.830 173.290 525.830 175.290 ;
        RECT 527.830 173.290 529.830 175.290 ;
        RECT 531.830 173.290 533.830 175.290 ;
        RECT 535.830 173.290 541.830 175.290 ;
        RECT 647.830 173.290 649.830 175.290 ;
        RECT 655.830 173.290 663.830 175.290 ;
        RECT 665.830 173.290 667.830 175.290 ;
        RECT 669.830 173.290 671.830 175.290 ;
        RECT 673.830 173.290 675.830 175.290 ;
        RECT 677.830 173.290 679.830 175.290 ;
        RECT 681.830 173.290 683.830 175.290 ;
        RECT 685.830 173.290 691.830 175.290 ;
        RECT 347.830 171.290 355.830 173.290 ;
        RECT 363.830 171.290 365.830 173.290 ;
        RECT 367.830 171.290 369.830 173.290 ;
        RECT 371.830 171.290 373.830 173.290 ;
        RECT 375.830 171.290 377.830 173.290 ;
        RECT 379.830 171.290 389.830 173.290 ;
        RECT 497.830 171.290 505.830 173.290 ;
        RECT 513.830 171.290 515.830 173.290 ;
        RECT 517.830 171.290 519.830 173.290 ;
        RECT 521.830 171.290 523.830 173.290 ;
        RECT 525.830 171.290 527.830 173.290 ;
        RECT 529.830 171.290 539.830 173.290 ;
        RECT 647.830 171.290 655.830 173.290 ;
        RECT 663.830 171.290 665.830 173.290 ;
        RECT 667.830 171.290 669.830 173.290 ;
        RECT 671.830 171.290 673.830 173.290 ;
        RECT 675.830 171.290 677.830 173.290 ;
        RECT 679.830 171.290 689.830 173.290 ;
        RECT 353.830 169.290 371.830 171.290 ;
        RECT 373.830 169.290 387.830 171.290 ;
        RECT 503.830 169.290 521.830 171.290 ;
        RECT 523.830 169.290 537.830 171.290 ;
        RECT 653.830 169.290 671.830 171.290 ;
        RECT 673.830 169.290 687.830 171.290 ;
        RECT 369.830 167.290 375.830 169.290 ;
        RECT 519.830 167.290 525.830 169.290 ;
        RECT 669.830 167.290 675.830 169.290 ;
        RECT 369.830 139.290 375.830 141.290 ;
        RECT 369.830 137.290 371.830 139.290 ;
        RECT 367.830 135.290 371.830 137.290 ;
        RECT 373.830 137.290 375.830 139.290 ;
        RECT 519.830 139.290 525.830 141.290 ;
        RECT 519.830 137.290 521.830 139.290 ;
        RECT 373.830 135.290 377.830 137.290 ;
        RECT 367.830 131.290 369.830 135.290 ;
        RECT 365.830 129.290 369.830 131.290 ;
        RECT 375.830 131.290 377.830 135.290 ;
        RECT 517.830 135.290 521.830 137.290 ;
        RECT 523.830 137.290 525.830 139.290 ;
        RECT 669.830 139.290 675.830 141.290 ;
        RECT 669.830 137.290 671.830 139.290 ;
        RECT 523.830 135.290 527.830 137.290 ;
        RECT 517.830 131.290 519.830 135.290 ;
        RECT 375.830 129.290 379.830 131.290 ;
        RECT 365.830 125.290 367.830 129.290 ;
        RECT 363.830 123.290 367.830 125.290 ;
        RECT 369.830 123.290 373.830 127.290 ;
        RECT 377.830 125.290 379.830 129.290 ;
        RECT 515.830 129.290 519.830 131.290 ;
        RECT 525.830 131.290 527.830 135.290 ;
        RECT 667.830 135.290 671.830 137.290 ;
        RECT 673.830 137.290 675.830 139.290 ;
        RECT 673.830 135.290 677.830 137.290 ;
        RECT 667.830 131.290 669.830 135.290 ;
        RECT 525.830 129.290 529.830 131.290 ;
        RECT 515.830 125.290 517.830 129.290 ;
        RECT 377.830 123.290 381.830 125.290 ;
        RECT 363.830 119.290 365.830 123.290 ;
        RECT 361.830 117.290 365.830 119.290 ;
        RECT 367.830 121.290 373.830 123.290 ;
        RECT 379.830 121.290 381.830 123.290 ;
        RECT 513.830 123.290 517.830 125.290 ;
        RECT 519.830 123.290 523.830 127.290 ;
        RECT 527.830 125.290 529.830 129.290 ;
        RECT 665.830 129.290 669.830 131.290 ;
        RECT 675.830 131.290 677.830 135.290 ;
        RECT 675.830 129.290 679.830 131.290 ;
        RECT 665.830 125.290 667.830 129.290 ;
        RECT 527.830 123.290 531.830 125.290 ;
        RECT 367.830 119.290 375.830 121.290 ;
        RECT 379.830 119.290 383.830 121.290 ;
        RECT 513.830 119.290 515.830 123.290 ;
        RECT 367.830 117.290 377.830 119.290 ;
        RECT 361.830 115.290 363.830 117.290 ;
        RECT 359.830 113.290 363.830 115.290 ;
        RECT 365.830 113.290 373.830 117.290 ;
        RECT 359.830 109.290 361.830 113.290 ;
        RECT 357.830 107.290 361.830 109.290 ;
        RECT 363.830 109.290 373.830 113.290 ;
        RECT 375.830 113.290 379.830 117.290 ;
        RECT 381.830 115.290 383.830 119.290 ;
        RECT 511.830 117.290 515.830 119.290 ;
        RECT 517.830 121.290 523.830 123.290 ;
        RECT 529.830 121.290 531.830 123.290 ;
        RECT 663.830 123.290 667.830 125.290 ;
        RECT 669.830 123.290 673.830 127.290 ;
        RECT 677.830 125.290 679.830 129.290 ;
        RECT 677.830 123.290 681.830 125.290 ;
        RECT 517.830 119.290 525.830 121.290 ;
        RECT 529.830 119.290 533.830 121.290 ;
        RECT 663.830 119.290 665.830 123.290 ;
        RECT 517.830 117.290 527.830 119.290 ;
        RECT 511.830 115.290 513.830 117.290 ;
        RECT 381.830 113.290 385.830 115.290 ;
        RECT 375.830 109.290 381.830 113.290 ;
        RECT 363.830 107.290 375.830 109.290 ;
        RECT 357.830 105.290 359.830 107.290 ;
        RECT 351.830 103.290 359.830 105.290 ;
        RECT 361.830 103.290 375.830 107.290 ;
        RECT 377.830 107.290 381.830 109.290 ;
        RECT 383.830 109.290 385.830 113.290 ;
        RECT 509.830 113.290 513.830 115.290 ;
        RECT 515.830 113.290 523.830 117.290 ;
        RECT 509.830 109.290 511.830 113.290 ;
        RECT 383.830 107.290 387.830 109.290 ;
        RECT 377.830 105.290 383.830 107.290 ;
        RECT 377.830 103.290 379.830 105.290 ;
        RECT 385.830 103.290 387.830 107.290 ;
        RECT 507.830 107.290 511.830 109.290 ;
        RECT 513.830 109.290 523.830 113.290 ;
        RECT 525.830 113.290 529.830 117.290 ;
        RECT 531.830 115.290 533.830 119.290 ;
        RECT 661.830 117.290 665.830 119.290 ;
        RECT 667.830 121.290 673.830 123.290 ;
        RECT 679.830 121.290 681.830 123.290 ;
        RECT 667.830 119.290 675.830 121.290 ;
        RECT 679.830 119.290 683.830 121.290 ;
        RECT 667.830 117.290 677.830 119.290 ;
        RECT 661.830 115.290 663.830 117.290 ;
        RECT 531.830 113.290 535.830 115.290 ;
        RECT 525.830 109.290 531.830 113.290 ;
        RECT 513.830 107.290 525.830 109.290 ;
        RECT 507.830 105.290 509.830 107.290 ;
        RECT 501.830 103.290 509.830 105.290 ;
        RECT 511.830 103.290 525.830 107.290 ;
        RECT 527.830 107.290 531.830 109.290 ;
        RECT 533.830 109.290 535.830 113.290 ;
        RECT 659.830 113.290 663.830 115.290 ;
        RECT 665.830 113.290 673.830 117.290 ;
        RECT 659.830 109.290 661.830 113.290 ;
        RECT 533.830 107.290 537.830 109.290 ;
        RECT 527.830 105.290 533.830 107.290 ;
        RECT 527.830 103.290 529.830 105.290 ;
        RECT 535.830 103.290 537.830 107.290 ;
        RECT 657.830 107.290 661.830 109.290 ;
        RECT 663.830 109.290 673.830 113.290 ;
        RECT 675.830 113.290 679.830 117.290 ;
        RECT 681.830 115.290 683.830 119.290 ;
        RECT 681.830 113.290 685.830 115.290 ;
        RECT 675.830 109.290 681.830 113.290 ;
        RECT 663.830 107.290 675.830 109.290 ;
        RECT 657.830 105.290 659.830 107.290 ;
        RECT 651.830 103.290 659.830 105.290 ;
        RECT 661.830 103.290 675.830 107.290 ;
        RECT 677.830 107.290 681.830 109.290 ;
        RECT 683.830 109.290 685.830 113.290 ;
        RECT 683.830 107.290 687.830 109.290 ;
        RECT 677.830 105.290 683.830 107.290 ;
        RECT 677.830 103.290 679.830 105.290 ;
        RECT 685.830 103.290 687.830 107.290 ;
        RECT 341.830 101.290 353.830 103.290 ;
        RECT 361.830 101.290 377.830 103.290 ;
        RECT 379.830 101.290 383.830 103.290 ;
        RECT 385.830 101.290 395.830 103.290 ;
        RECT 491.830 101.290 503.830 103.290 ;
        RECT 511.830 101.290 527.830 103.290 ;
        RECT 529.830 101.290 533.830 103.290 ;
        RECT 535.830 101.290 545.830 103.290 ;
        RECT 641.830 101.290 653.830 103.290 ;
        RECT 661.830 101.290 677.830 103.290 ;
        RECT 679.830 101.290 683.830 103.290 ;
        RECT 685.830 101.290 695.830 103.290 ;
        RECT 335.830 99.290 343.830 101.290 ;
        RECT 353.830 99.290 357.830 101.290 ;
        RECT 335.830 95.290 337.830 99.290 ;
        RECT 343.830 97.290 357.830 99.290 ;
        RECT 359.830 97.290 385.830 101.290 ;
        RECT 393.830 99.290 403.830 101.290 ;
        RECT 485.830 99.290 493.830 101.290 ;
        RECT 503.830 99.290 507.830 101.290 ;
        RECT 387.830 97.290 389.830 99.290 ;
        RECT 401.830 97.290 411.830 99.290 ;
        RECT 343.830 95.290 359.830 97.290 ;
        RECT 369.830 95.290 381.830 97.290 ;
        RECT 385.830 95.290 393.830 97.290 ;
        RECT 409.830 95.290 415.830 97.290 ;
        RECT 335.830 93.290 343.830 95.290 ;
        RECT 353.830 93.290 369.830 95.290 ;
        RECT 381.830 93.290 399.830 95.290 ;
        RECT 413.830 93.290 415.830 95.290 ;
        RECT 485.830 95.290 487.830 99.290 ;
        RECT 493.830 97.290 507.830 99.290 ;
        RECT 509.830 97.290 535.830 101.290 ;
        RECT 543.830 99.290 553.830 101.290 ;
        RECT 635.830 99.290 643.830 101.290 ;
        RECT 653.830 99.290 657.830 101.290 ;
        RECT 537.830 97.290 539.830 99.290 ;
        RECT 551.830 97.290 561.830 99.290 ;
        RECT 493.830 95.290 509.830 97.290 ;
        RECT 519.830 95.290 531.830 97.290 ;
        RECT 535.830 95.290 543.830 97.290 ;
        RECT 559.830 95.290 565.830 97.290 ;
        RECT 485.830 93.290 493.830 95.290 ;
        RECT 503.830 93.290 519.830 95.290 ;
        RECT 531.830 93.290 549.830 95.290 ;
        RECT 563.830 93.290 565.830 95.290 ;
        RECT 635.830 95.290 637.830 99.290 ;
        RECT 643.830 97.290 657.830 99.290 ;
        RECT 659.830 97.290 685.830 101.290 ;
        RECT 693.830 99.290 703.830 101.290 ;
        RECT 687.830 97.290 689.830 99.290 ;
        RECT 701.830 97.290 711.830 99.290 ;
        RECT 643.830 95.290 659.830 97.290 ;
        RECT 669.830 95.290 681.830 97.290 ;
        RECT 685.830 95.290 693.830 97.290 ;
        RECT 709.830 95.290 715.830 97.290 ;
        RECT 635.830 93.290 643.830 95.290 ;
        RECT 653.830 93.290 669.830 95.290 ;
        RECT 681.830 93.290 699.830 95.290 ;
        RECT 713.830 93.290 715.830 95.290 ;
        RECT 341.830 91.290 353.830 93.290 ;
        RECT 363.830 91.290 403.830 93.290 ;
        RECT 411.830 91.290 415.830 93.290 ;
        RECT 491.830 91.290 503.830 93.290 ;
        RECT 513.830 91.290 553.830 93.290 ;
        RECT 561.830 91.290 565.830 93.290 ;
        RECT 641.830 91.290 653.830 93.290 ;
        RECT 663.830 91.290 703.830 93.290 ;
        RECT 711.830 91.290 715.830 93.290 ;
        RECT 351.830 89.290 363.830 91.290 ;
        RECT 373.830 89.290 401.830 91.290 ;
        RECT 409.830 89.290 413.830 91.290 ;
        RECT 501.830 89.290 513.830 91.290 ;
        RECT 523.830 89.290 551.830 91.290 ;
        RECT 559.830 89.290 563.830 91.290 ;
        RECT 651.830 89.290 663.830 91.290 ;
        RECT 673.830 89.290 701.830 91.290 ;
        RECT 709.830 89.290 713.830 91.290 ;
        RECT 353.830 87.290 355.830 89.290 ;
        RECT 351.830 85.290 355.830 87.290 ;
        RECT 357.830 87.290 373.830 89.290 ;
        RECT 383.830 87.290 393.830 89.290 ;
        RECT 401.830 87.290 411.830 89.290 ;
        RECT 503.830 87.290 505.830 89.290 ;
        RECT 357.830 85.290 383.830 87.290 ;
        RECT 393.830 85.290 403.830 87.290 ;
        RECT 501.830 85.290 505.830 87.290 ;
        RECT 507.830 87.290 523.830 89.290 ;
        RECT 533.830 87.290 543.830 89.290 ;
        RECT 551.830 87.290 561.830 89.290 ;
        RECT 653.830 87.290 655.830 89.290 ;
        RECT 507.830 85.290 533.830 87.290 ;
        RECT 543.830 85.290 553.830 87.290 ;
        RECT 651.830 85.290 655.830 87.290 ;
        RECT 657.830 87.290 673.830 89.290 ;
        RECT 683.830 87.290 693.830 89.290 ;
        RECT 701.830 87.290 711.830 89.290 ;
        RECT 657.830 85.290 683.830 87.290 ;
        RECT 693.830 85.290 703.830 87.290 ;
        RECT 351.830 79.290 353.830 85.290 ;
        RECT 355.830 83.290 373.830 85.290 ;
        RECT 383.830 83.290 395.830 85.290 ;
        RECT 355.830 81.290 371.830 83.290 ;
        RECT 357.830 79.290 371.830 81.290 ;
        RECT 373.830 81.290 377.830 83.290 ;
        RECT 381.830 81.290 383.830 83.290 ;
        RECT 387.830 81.290 389.830 83.290 ;
        RECT 393.830 81.290 395.830 83.290 ;
        RECT 403.830 81.290 409.830 83.290 ;
        RECT 373.830 79.290 375.830 81.290 ;
        RECT 387.830 79.290 395.830 81.290 ;
        RECT 401.830 79.290 405.830 81.290 ;
        RECT 407.830 79.290 409.830 81.290 ;
        RECT 501.830 79.290 503.830 85.290 ;
        RECT 505.830 83.290 523.830 85.290 ;
        RECT 533.830 83.290 545.830 85.290 ;
        RECT 505.830 81.290 521.830 83.290 ;
        RECT 507.830 79.290 521.830 81.290 ;
        RECT 523.830 81.290 527.830 83.290 ;
        RECT 531.830 81.290 533.830 83.290 ;
        RECT 537.830 81.290 539.830 83.290 ;
        RECT 543.830 81.290 545.830 83.290 ;
        RECT 553.830 81.290 559.830 83.290 ;
        RECT 523.830 79.290 525.830 81.290 ;
        RECT 537.830 79.290 545.830 81.290 ;
        RECT 551.830 79.290 555.830 81.290 ;
        RECT 557.830 79.290 559.830 81.290 ;
        RECT 651.830 79.290 653.830 85.290 ;
        RECT 655.830 83.290 673.830 85.290 ;
        RECT 683.830 83.290 695.830 85.290 ;
        RECT 655.830 81.290 671.830 83.290 ;
        RECT 657.830 79.290 671.830 81.290 ;
        RECT 673.830 81.290 677.830 83.290 ;
        RECT 681.830 81.290 683.830 83.290 ;
        RECT 687.830 81.290 689.830 83.290 ;
        RECT 693.830 81.290 695.830 83.290 ;
        RECT 703.830 81.290 709.830 83.290 ;
        RECT 673.830 79.290 675.830 81.290 ;
        RECT 687.830 79.290 695.830 81.290 ;
        RECT 701.830 79.290 705.830 81.290 ;
        RECT 707.830 79.290 709.830 81.290 ;
        RECT 349.830 77.290 355.830 79.290 ;
        RECT 347.830 75.290 351.830 77.290 ;
        RECT 353.830 75.290 359.830 77.290 ;
        RECT 361.830 75.290 371.830 79.290 ;
        RECT 375.830 77.290 377.830 79.290 ;
        RECT 387.830 77.290 391.830 79.290 ;
        RECT 397.830 77.290 403.830 79.290 ;
        RECT 405.830 77.290 409.830 79.290 ;
        RECT 499.830 77.290 505.830 79.290 ;
        RECT 385.830 75.290 391.830 77.290 ;
        RECT 393.830 75.290 399.830 77.290 ;
        RECT 345.830 73.290 349.830 75.290 ;
        RECT 351.830 73.290 361.830 75.290 ;
        RECT 365.830 73.290 373.830 75.290 ;
        RECT 379.830 73.290 395.830 75.290 ;
        RECT 399.830 73.290 403.830 75.290 ;
        RECT 5.000 60.000 25.000 70.000 ;
        RECT 345.830 67.290 347.830 73.290 ;
        RECT 343.830 65.290 347.830 67.290 ;
        RECT 349.830 71.290 363.830 73.290 ;
        RECT 367.830 71.290 373.830 73.290 ;
        RECT 383.830 71.290 391.830 73.290 ;
        RECT 395.830 71.290 405.830 73.290 ;
        RECT 407.830 71.290 409.830 77.290 ;
        RECT 497.830 75.290 501.830 77.290 ;
        RECT 503.830 75.290 509.830 77.290 ;
        RECT 511.830 75.290 521.830 79.290 ;
        RECT 525.830 77.290 527.830 79.290 ;
        RECT 537.830 77.290 541.830 79.290 ;
        RECT 547.830 77.290 553.830 79.290 ;
        RECT 555.830 77.290 559.830 79.290 ;
        RECT 649.830 77.290 655.830 79.290 ;
        RECT 535.830 75.290 541.830 77.290 ;
        RECT 543.830 75.290 549.830 77.290 ;
        RECT 349.830 69.290 367.830 71.290 ;
        RECT 369.830 69.290 373.830 71.290 ;
        RECT 381.830 69.290 387.830 71.290 ;
        RECT 391.830 69.290 401.830 71.290 ;
        RECT 405.830 69.290 409.830 71.290 ;
        RECT 495.830 73.290 499.830 75.290 ;
        RECT 501.830 73.290 511.830 75.290 ;
        RECT 515.830 73.290 523.830 75.290 ;
        RECT 529.830 73.290 545.830 75.290 ;
        RECT 549.830 73.290 553.830 75.290 ;
        RECT 349.830 67.290 369.830 69.290 ;
        RECT 377.830 67.290 383.830 69.290 ;
        RECT 387.830 67.290 399.830 69.290 ;
        RECT 349.830 65.290 389.830 67.290 ;
        RECT 397.830 65.290 399.830 67.290 ;
        RECT 401.830 67.290 407.830 69.290 ;
        RECT 495.830 67.290 497.830 73.290 ;
        RECT 401.830 65.290 403.830 67.290 ;
        RECT 343.830 45.290 345.830 65.290 ;
        RECT 347.830 63.290 363.830 65.290 ;
        RECT 365.830 63.290 367.830 65.290 ;
        RECT 371.830 63.290 383.830 65.290 ;
        RECT 347.830 61.290 361.830 63.290 ;
        RECT 363.830 61.290 365.830 63.290 ;
        RECT 367.830 61.290 371.830 63.290 ;
        RECT 377.830 61.290 381.830 63.290 ;
        RECT 383.830 61.290 385.830 63.290 ;
        RECT 399.830 61.290 403.830 65.290 ;
        RECT 347.830 59.290 363.830 61.290 ;
        RECT 365.830 59.290 367.830 61.290 ;
        RECT 347.830 57.290 361.830 59.290 ;
        RECT 363.830 57.290 367.830 59.290 ;
        RECT 371.830 59.290 381.830 61.290 ;
        RECT 385.830 59.290 403.830 61.290 ;
        RECT 493.830 65.290 497.830 67.290 ;
        RECT 499.830 71.290 513.830 73.290 ;
        RECT 517.830 71.290 523.830 73.290 ;
        RECT 533.830 71.290 541.830 73.290 ;
        RECT 545.830 71.290 555.830 73.290 ;
        RECT 557.830 71.290 559.830 77.290 ;
        RECT 647.830 75.290 651.830 77.290 ;
        RECT 653.830 75.290 659.830 77.290 ;
        RECT 661.830 75.290 671.830 79.290 ;
        RECT 675.830 77.290 677.830 79.290 ;
        RECT 687.830 77.290 691.830 79.290 ;
        RECT 697.830 77.290 703.830 79.290 ;
        RECT 705.830 77.290 709.830 79.290 ;
        RECT 685.830 75.290 691.830 77.290 ;
        RECT 693.830 75.290 699.830 77.290 ;
        RECT 499.830 69.290 517.830 71.290 ;
        RECT 519.830 69.290 523.830 71.290 ;
        RECT 531.830 69.290 537.830 71.290 ;
        RECT 541.830 69.290 551.830 71.290 ;
        RECT 555.830 69.290 559.830 71.290 ;
        RECT 645.830 73.290 649.830 75.290 ;
        RECT 651.830 73.290 661.830 75.290 ;
        RECT 665.830 73.290 673.830 75.290 ;
        RECT 679.830 73.290 695.830 75.290 ;
        RECT 699.830 73.290 703.830 75.290 ;
        RECT 499.830 67.290 519.830 69.290 ;
        RECT 527.830 67.290 533.830 69.290 ;
        RECT 537.830 67.290 549.830 69.290 ;
        RECT 499.830 65.290 539.830 67.290 ;
        RECT 547.830 65.290 549.830 67.290 ;
        RECT 551.830 67.290 557.830 69.290 ;
        RECT 645.830 67.290 647.830 73.290 ;
        RECT 551.830 65.290 553.830 67.290 ;
        RECT 371.830 57.290 373.830 59.290 ;
        RECT 379.830 57.290 383.830 59.290 ;
        RECT 387.830 57.290 389.830 59.290 ;
        RECT 401.830 57.290 405.830 59.290 ;
        RECT 347.830 55.290 363.830 57.290 ;
        RECT 365.830 55.290 367.830 57.290 ;
        RECT 373.830 55.290 377.830 57.290 ;
        RECT 347.830 53.290 365.830 55.290 ;
        RECT 367.830 53.290 369.830 55.290 ;
        RECT 375.830 53.290 377.830 55.290 ;
        RECT 379.830 55.290 381.830 57.290 ;
        RECT 379.830 53.290 383.830 55.290 ;
        RECT 385.830 53.290 387.830 57.290 ;
        RECT 403.830 55.290 407.830 57.290 ;
        RECT 399.830 53.290 403.830 55.290 ;
        RECT 347.830 51.290 363.830 53.290 ;
        RECT 369.830 51.290 371.830 53.290 ;
        RECT 377.830 51.290 385.830 53.290 ;
        RECT 387.830 51.290 391.830 53.290 ;
        RECT 395.830 51.290 401.830 53.290 ;
        RECT 405.830 51.290 407.830 55.290 ;
        RECT 347.830 49.290 365.830 51.290 ;
        RECT 371.830 49.290 373.830 51.290 ;
        RECT 381.830 49.290 387.830 51.290 ;
        RECT 391.830 49.290 395.830 51.290 ;
        RECT 401.830 49.290 407.830 51.290 ;
        RECT 347.830 47.290 363.830 49.290 ;
        RECT 373.830 47.290 375.830 49.290 ;
        RECT 383.830 47.290 391.830 49.290 ;
        RECT 395.830 47.290 403.830 49.290 ;
        RECT 347.830 45.290 361.830 47.290 ;
        RECT 363.830 45.290 365.830 47.290 ;
        RECT 375.830 45.290 379.830 47.290 ;
        RECT 389.830 45.290 397.830 47.290 ;
        RECT 493.830 45.290 495.830 65.290 ;
        RECT 497.830 63.290 513.830 65.290 ;
        RECT 515.830 63.290 517.830 65.290 ;
        RECT 521.830 63.290 533.830 65.290 ;
        RECT 497.830 61.290 511.830 63.290 ;
        RECT 513.830 61.290 515.830 63.290 ;
        RECT 517.830 61.290 521.830 63.290 ;
        RECT 527.830 61.290 531.830 63.290 ;
        RECT 533.830 61.290 535.830 63.290 ;
        RECT 549.830 61.290 553.830 65.290 ;
        RECT 497.830 59.290 513.830 61.290 ;
        RECT 515.830 59.290 517.830 61.290 ;
        RECT 497.830 57.290 511.830 59.290 ;
        RECT 513.830 57.290 517.830 59.290 ;
        RECT 521.830 59.290 531.830 61.290 ;
        RECT 535.830 59.290 553.830 61.290 ;
        RECT 643.830 65.290 647.830 67.290 ;
        RECT 649.830 71.290 663.830 73.290 ;
        RECT 667.830 71.290 673.830 73.290 ;
        RECT 683.830 71.290 691.830 73.290 ;
        RECT 695.830 71.290 705.830 73.290 ;
        RECT 707.830 71.290 709.830 77.290 ;
        RECT 649.830 69.290 667.830 71.290 ;
        RECT 669.830 69.290 673.830 71.290 ;
        RECT 681.830 69.290 687.830 71.290 ;
        RECT 691.830 69.290 701.830 71.290 ;
        RECT 705.830 69.290 709.830 71.290 ;
        RECT 649.830 67.290 669.830 69.290 ;
        RECT 677.830 67.290 683.830 69.290 ;
        RECT 687.830 67.290 699.830 69.290 ;
        RECT 649.830 65.290 689.830 67.290 ;
        RECT 697.830 65.290 699.830 67.290 ;
        RECT 701.830 67.290 707.830 69.290 ;
        RECT 701.830 65.290 703.830 67.290 ;
        RECT 521.830 57.290 523.830 59.290 ;
        RECT 529.830 57.290 533.830 59.290 ;
        RECT 537.830 57.290 539.830 59.290 ;
        RECT 551.830 57.290 555.830 59.290 ;
        RECT 497.830 55.290 513.830 57.290 ;
        RECT 515.830 55.290 517.830 57.290 ;
        RECT 523.830 55.290 527.830 57.290 ;
        RECT 497.830 53.290 515.830 55.290 ;
        RECT 517.830 53.290 519.830 55.290 ;
        RECT 525.830 53.290 527.830 55.290 ;
        RECT 529.830 55.290 531.830 57.290 ;
        RECT 529.830 53.290 533.830 55.290 ;
        RECT 535.830 53.290 537.830 57.290 ;
        RECT 553.830 55.290 557.830 57.290 ;
        RECT 549.830 53.290 553.830 55.290 ;
        RECT 497.830 51.290 513.830 53.290 ;
        RECT 519.830 51.290 521.830 53.290 ;
        RECT 527.830 51.290 535.830 53.290 ;
        RECT 537.830 51.290 541.830 53.290 ;
        RECT 545.830 51.290 551.830 53.290 ;
        RECT 555.830 51.290 557.830 55.290 ;
        RECT 497.830 49.290 515.830 51.290 ;
        RECT 521.830 49.290 523.830 51.290 ;
        RECT 531.830 49.290 537.830 51.290 ;
        RECT 541.830 49.290 545.830 51.290 ;
        RECT 551.830 49.290 557.830 51.290 ;
        RECT 497.830 47.290 513.830 49.290 ;
        RECT 523.830 47.290 525.830 49.290 ;
        RECT 533.830 47.290 541.830 49.290 ;
        RECT 545.830 47.290 553.830 49.290 ;
        RECT 497.830 45.290 511.830 47.290 ;
        RECT 513.830 45.290 515.830 47.290 ;
        RECT 525.830 45.290 529.830 47.290 ;
        RECT 539.830 45.290 547.830 47.290 ;
        RECT 643.830 45.290 645.830 65.290 ;
        RECT 647.830 63.290 663.830 65.290 ;
        RECT 665.830 63.290 667.830 65.290 ;
        RECT 671.830 63.290 683.830 65.290 ;
        RECT 647.830 61.290 661.830 63.290 ;
        RECT 663.830 61.290 665.830 63.290 ;
        RECT 667.830 61.290 671.830 63.290 ;
        RECT 677.830 61.290 681.830 63.290 ;
        RECT 683.830 61.290 685.830 63.290 ;
        RECT 699.830 61.290 703.830 65.290 ;
        RECT 647.830 59.290 663.830 61.290 ;
        RECT 665.830 59.290 667.830 61.290 ;
        RECT 647.830 57.290 661.830 59.290 ;
        RECT 663.830 57.290 667.830 59.290 ;
        RECT 671.830 59.290 681.830 61.290 ;
        RECT 685.830 59.290 703.830 61.290 ;
        RECT 671.830 57.290 673.830 59.290 ;
        RECT 679.830 57.290 683.830 59.290 ;
        RECT 687.830 57.290 689.830 59.290 ;
        RECT 701.830 57.290 705.830 59.290 ;
        RECT 647.830 55.290 663.830 57.290 ;
        RECT 665.830 55.290 667.830 57.290 ;
        RECT 673.830 55.290 677.830 57.290 ;
        RECT 647.830 53.290 665.830 55.290 ;
        RECT 667.830 53.290 669.830 55.290 ;
        RECT 675.830 53.290 677.830 55.290 ;
        RECT 679.830 55.290 681.830 57.290 ;
        RECT 679.830 53.290 683.830 55.290 ;
        RECT 685.830 53.290 687.830 57.290 ;
        RECT 703.830 55.290 707.830 57.290 ;
        RECT 699.830 53.290 703.830 55.290 ;
        RECT 647.830 51.290 663.830 53.290 ;
        RECT 669.830 51.290 671.830 53.290 ;
        RECT 677.830 51.290 685.830 53.290 ;
        RECT 687.830 51.290 691.830 53.290 ;
        RECT 695.830 51.290 701.830 53.290 ;
        RECT 705.830 51.290 707.830 55.290 ;
        RECT 647.830 49.290 665.830 51.290 ;
        RECT 671.830 49.290 673.830 51.290 ;
        RECT 681.830 49.290 687.830 51.290 ;
        RECT 691.830 49.290 695.830 51.290 ;
        RECT 701.830 49.290 707.830 51.290 ;
        RECT 647.830 47.290 663.830 49.290 ;
        RECT 673.830 47.290 675.830 49.290 ;
        RECT 683.830 47.290 691.830 49.290 ;
        RECT 695.830 47.290 703.830 49.290 ;
        RECT 647.830 45.290 661.830 47.290 ;
        RECT 663.830 45.290 665.830 47.290 ;
        RECT 675.830 45.290 679.830 47.290 ;
        RECT 689.830 45.290 697.830 47.290 ;
        RECT 343.830 43.290 347.830 45.290 ;
        RECT 85.000 30.000 105.000 40.000 ;
        RECT 345.830 27.290 347.830 43.290 ;
        RECT 349.830 41.290 359.830 45.290 ;
        RECT 361.830 43.290 363.830 45.290 ;
        RECT 365.830 43.290 367.830 45.290 ;
        RECT 379.830 43.290 393.830 45.290 ;
        RECT 493.830 43.290 497.830 45.290 ;
        RECT 363.830 41.290 365.830 43.290 ;
        RECT 379.830 41.290 389.830 43.290 ;
        RECT 349.830 39.290 363.830 41.290 ;
        RECT 365.830 39.290 367.830 41.290 ;
        RECT 381.830 39.290 389.830 41.290 ;
        RECT 349.830 37.290 361.830 39.290 ;
        RECT 363.830 37.290 365.830 39.290 ;
        RECT 349.830 35.290 363.830 37.290 ;
        RECT 365.830 35.290 367.830 37.290 ;
        RECT 381.830 35.290 391.830 39.290 ;
        RECT 349.830 33.290 365.830 35.290 ;
        RECT 349.830 31.290 363.830 33.290 ;
        RECT 365.830 31.290 367.830 33.290 ;
        RECT 383.830 31.290 391.830 35.290 ;
        RECT 349.830 29.290 365.830 31.290 ;
        RECT 349.830 27.290 363.830 29.290 ;
        RECT 365.830 27.290 367.830 29.290 ;
        RECT 385.830 27.290 391.830 31.290 ;
        RECT 345.830 25.290 349.830 27.290 ;
        RECT 351.830 25.290 365.830 27.290 ;
        RECT 383.830 25.290 385.830 27.290 ;
        RECT 389.830 25.290 391.830 27.290 ;
        RECT 495.830 27.290 497.830 43.290 ;
        RECT 499.830 41.290 509.830 45.290 ;
        RECT 511.830 43.290 513.830 45.290 ;
        RECT 515.830 43.290 517.830 45.290 ;
        RECT 529.830 43.290 543.830 45.290 ;
        RECT 643.830 43.290 647.830 45.290 ;
        RECT 513.830 41.290 515.830 43.290 ;
        RECT 529.830 41.290 539.830 43.290 ;
        RECT 499.830 39.290 513.830 41.290 ;
        RECT 515.830 39.290 517.830 41.290 ;
        RECT 531.830 39.290 539.830 41.290 ;
        RECT 499.830 37.290 511.830 39.290 ;
        RECT 513.830 37.290 515.830 39.290 ;
        RECT 499.830 35.290 513.830 37.290 ;
        RECT 515.830 35.290 517.830 37.290 ;
        RECT 531.830 35.290 541.830 39.290 ;
        RECT 499.830 33.290 515.830 35.290 ;
        RECT 499.830 31.290 513.830 33.290 ;
        RECT 515.830 31.290 517.830 33.290 ;
        RECT 533.830 31.290 541.830 35.290 ;
        RECT 499.830 29.290 515.830 31.290 ;
        RECT 499.830 27.290 513.830 29.290 ;
        RECT 515.830 27.290 517.830 29.290 ;
        RECT 535.830 27.290 541.830 31.290 ;
        RECT 495.830 25.290 499.830 27.290 ;
        RECT 501.830 25.290 515.830 27.290 ;
        RECT 533.830 25.290 535.830 27.290 ;
        RECT 539.830 25.290 541.830 27.290 ;
        RECT 645.830 27.290 647.830 43.290 ;
        RECT 649.830 41.290 659.830 45.290 ;
        RECT 661.830 43.290 663.830 45.290 ;
        RECT 665.830 43.290 667.830 45.290 ;
        RECT 679.830 43.290 693.830 45.290 ;
        RECT 663.830 41.290 665.830 43.290 ;
        RECT 679.830 41.290 689.830 43.290 ;
        RECT 649.830 39.290 663.830 41.290 ;
        RECT 665.830 39.290 667.830 41.290 ;
        RECT 681.830 39.290 689.830 41.290 ;
        RECT 649.830 37.290 661.830 39.290 ;
        RECT 663.830 37.290 665.830 39.290 ;
        RECT 649.830 35.290 663.830 37.290 ;
        RECT 665.830 35.290 667.830 37.290 ;
        RECT 681.830 35.290 691.830 39.290 ;
        RECT 649.830 33.290 665.830 35.290 ;
        RECT 649.830 31.290 663.830 33.290 ;
        RECT 665.830 31.290 667.830 33.290 ;
        RECT 683.830 31.290 691.830 35.290 ;
        RECT 649.830 29.290 665.830 31.290 ;
        RECT 649.830 27.290 663.830 29.290 ;
        RECT 665.830 27.290 667.830 29.290 ;
        RECT 685.830 27.290 691.830 31.290 ;
        RECT 645.830 25.290 649.830 27.290 ;
        RECT 651.830 25.290 665.830 27.290 ;
        RECT 683.830 25.290 685.830 27.290 ;
        RECT 689.830 25.290 691.830 27.290 ;
        RECT 85.000 5.000 105.000 25.000 ;
        RECT 347.830 23.290 349.830 25.290 ;
        RECT 355.830 23.290 363.830 25.290 ;
        RECT 365.830 23.290 367.830 25.290 ;
        RECT 369.830 23.290 371.830 25.290 ;
        RECT 373.830 23.290 375.830 25.290 ;
        RECT 377.830 23.290 379.830 25.290 ;
        RECT 381.830 23.290 383.830 25.290 ;
        RECT 385.830 23.290 391.830 25.290 ;
        RECT 497.830 23.290 499.830 25.290 ;
        RECT 505.830 23.290 513.830 25.290 ;
        RECT 515.830 23.290 517.830 25.290 ;
        RECT 519.830 23.290 521.830 25.290 ;
        RECT 523.830 23.290 525.830 25.290 ;
        RECT 527.830 23.290 529.830 25.290 ;
        RECT 531.830 23.290 533.830 25.290 ;
        RECT 535.830 23.290 541.830 25.290 ;
        RECT 647.830 23.290 649.830 25.290 ;
        RECT 655.830 23.290 663.830 25.290 ;
        RECT 665.830 23.290 667.830 25.290 ;
        RECT 669.830 23.290 671.830 25.290 ;
        RECT 673.830 23.290 675.830 25.290 ;
        RECT 677.830 23.290 679.830 25.290 ;
        RECT 681.830 23.290 683.830 25.290 ;
        RECT 685.830 23.290 691.830 25.290 ;
        RECT 347.830 21.290 355.830 23.290 ;
        RECT 363.830 21.290 365.830 23.290 ;
        RECT 367.830 21.290 369.830 23.290 ;
        RECT 371.830 21.290 373.830 23.290 ;
        RECT 375.830 21.290 377.830 23.290 ;
        RECT 379.830 21.290 389.830 23.290 ;
        RECT 497.830 21.290 505.830 23.290 ;
        RECT 513.830 21.290 515.830 23.290 ;
        RECT 517.830 21.290 519.830 23.290 ;
        RECT 521.830 21.290 523.830 23.290 ;
        RECT 525.830 21.290 527.830 23.290 ;
        RECT 529.830 21.290 539.830 23.290 ;
        RECT 647.830 21.290 655.830 23.290 ;
        RECT 663.830 21.290 665.830 23.290 ;
        RECT 667.830 21.290 669.830 23.290 ;
        RECT 671.830 21.290 673.830 23.290 ;
        RECT 675.830 21.290 677.830 23.290 ;
        RECT 679.830 21.290 689.830 23.290 ;
        RECT 353.830 19.290 371.830 21.290 ;
        RECT 373.830 19.290 387.830 21.290 ;
        RECT 503.830 19.290 521.830 21.290 ;
        RECT 523.830 19.290 537.830 21.290 ;
        RECT 653.830 19.290 671.830 21.290 ;
        RECT 673.830 19.290 687.830 21.290 ;
        RECT 369.830 17.290 375.830 19.290 ;
        RECT 519.830 17.290 525.830 19.290 ;
        RECT 669.830 17.290 675.830 19.290 ;
        RECT 749.000 0.000 749.800 300.000 ;
  END
END Art
END LIBRARY

