* NGSPICE file created from ExperiarCore.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

.subckt ExperiarCore addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] addr0[8] addr1[0] addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6]
+ addr1[7] addr1[8] clk0 clk1 coreIndex[0] coreIndex[1] coreIndex[2] coreIndex[3]
+ coreIndex[4] coreIndex[5] coreIndex[6] coreIndex[7] core_wb_ack_i core_wb_adr_o[0]
+ core_wb_adr_o[10] core_wb_adr_o[11] core_wb_adr_o[12] core_wb_adr_o[13] core_wb_adr_o[14]
+ core_wb_adr_o[15] core_wb_adr_o[16] core_wb_adr_o[17] core_wb_adr_o[18] core_wb_adr_o[19]
+ core_wb_adr_o[1] core_wb_adr_o[20] core_wb_adr_o[21] core_wb_adr_o[22] core_wb_adr_o[23]
+ core_wb_adr_o[24] core_wb_adr_o[25] core_wb_adr_o[26] core_wb_adr_o[27] core_wb_adr_o[2]
+ core_wb_adr_o[3] core_wb_adr_o[4] core_wb_adr_o[5] core_wb_adr_o[6] core_wb_adr_o[7]
+ core_wb_adr_o[8] core_wb_adr_o[9] core_wb_cyc_o core_wb_data_i[0] core_wb_data_i[10]
+ core_wb_data_i[11] core_wb_data_i[12] core_wb_data_i[13] core_wb_data_i[14] core_wb_data_i[15]
+ core_wb_data_i[16] core_wb_data_i[17] core_wb_data_i[18] core_wb_data_i[19] core_wb_data_i[1]
+ core_wb_data_i[20] core_wb_data_i[21] core_wb_data_i[22] core_wb_data_i[23] core_wb_data_i[24]
+ core_wb_data_i[25] core_wb_data_i[26] core_wb_data_i[27] core_wb_data_i[28] core_wb_data_i[29]
+ core_wb_data_i[2] core_wb_data_i[30] core_wb_data_i[31] core_wb_data_i[3] core_wb_data_i[4]
+ core_wb_data_i[5] core_wb_data_i[6] core_wb_data_i[7] core_wb_data_i[8] core_wb_data_i[9]
+ core_wb_data_o[0] core_wb_data_o[10] core_wb_data_o[11] core_wb_data_o[12] core_wb_data_o[13]
+ core_wb_data_o[14] core_wb_data_o[15] core_wb_data_o[16] core_wb_data_o[17] core_wb_data_o[18]
+ core_wb_data_o[19] core_wb_data_o[1] core_wb_data_o[20] core_wb_data_o[21] core_wb_data_o[22]
+ core_wb_data_o[23] core_wb_data_o[24] core_wb_data_o[25] core_wb_data_o[26] core_wb_data_o[27]
+ core_wb_data_o[28] core_wb_data_o[29] core_wb_data_o[2] core_wb_data_o[30] core_wb_data_o[31]
+ core_wb_data_o[3] core_wb_data_o[4] core_wb_data_o[5] core_wb_data_o[6] core_wb_data_o[7]
+ core_wb_data_o[8] core_wb_data_o[9] core_wb_error_i core_wb_sel_o[0] core_wb_sel_o[1]
+ core_wb_sel_o[2] core_wb_sel_o[3] core_wb_stall_i core_wb_stb_o core_wb_we_o csb0[0]
+ csb0[1] csb1[0] csb1[1] din0[0] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[1] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[2] din0[30] din0[31]
+ din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] dout0[0] dout0[10] dout0[11]
+ dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19]
+ dout0[1] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[2] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34] dout0[35]
+ dout0[36] dout0[37] dout0[38] dout0[39] dout0[3] dout0[40] dout0[41] dout0[42] dout0[43]
+ dout0[44] dout0[45] dout0[46] dout0[47] dout0[48] dout0[49] dout0[4] dout0[50] dout0[51]
+ dout0[52] dout0[53] dout0[54] dout0[55] dout0[56] dout0[57] dout0[58] dout0[59]
+ dout0[5] dout0[60] dout0[61] dout0[62] dout0[63] dout0[6] dout0[7] dout0[8] dout0[9]
+ dout1[0] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16] dout1[17]
+ dout1[18] dout1[19] dout1[1] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24] dout1[25]
+ dout1[26] dout1[27] dout1[28] dout1[29] dout1[2] dout1[30] dout1[31] dout1[32] dout1[33]
+ dout1[34] dout1[35] dout1[36] dout1[37] dout1[38] dout1[39] dout1[3] dout1[40] dout1[41]
+ dout1[42] dout1[43] dout1[44] dout1[45] dout1[46] dout1[47] dout1[48] dout1[49]
+ dout1[4] dout1[50] dout1[51] dout1[52] dout1[53] dout1[54] dout1[55] dout1[56] dout1[57]
+ dout1[58] dout1[59] dout1[5] dout1[60] dout1[61] dout1[62] dout1[63] dout1[6] dout1[7]
+ dout1[8] dout1[9] irq[0] irq[10] irq[11] irq[12] irq[13] irq[14] irq[15] irq[1]
+ irq[2] irq[3] irq[4] irq[5] irq[6] irq[7] irq[8] irq[9] jtag_tck jtag_tdi jtag_tdo
+ jtag_tms localMemory_wb_ack_o localMemory_wb_adr_i[0] localMemory_wb_adr_i[10] localMemory_wb_adr_i[11]
+ localMemory_wb_adr_i[12] localMemory_wb_adr_i[13] localMemory_wb_adr_i[14] localMemory_wb_adr_i[15]
+ localMemory_wb_adr_i[16] localMemory_wb_adr_i[17] localMemory_wb_adr_i[18] localMemory_wb_adr_i[19]
+ localMemory_wb_adr_i[1] localMemory_wb_adr_i[20] localMemory_wb_adr_i[21] localMemory_wb_adr_i[22]
+ localMemory_wb_adr_i[23] localMemory_wb_adr_i[2] localMemory_wb_adr_i[3] localMemory_wb_adr_i[4]
+ localMemory_wb_adr_i[5] localMemory_wb_adr_i[6] localMemory_wb_adr_i[7] localMemory_wb_adr_i[8]
+ localMemory_wb_adr_i[9] localMemory_wb_cyc_i localMemory_wb_data_i[0] localMemory_wb_data_i[10]
+ localMemory_wb_data_i[11] localMemory_wb_data_i[12] localMemory_wb_data_i[13] localMemory_wb_data_i[14]
+ localMemory_wb_data_i[15] localMemory_wb_data_i[16] localMemory_wb_data_i[17] localMemory_wb_data_i[18]
+ localMemory_wb_data_i[19] localMemory_wb_data_i[1] localMemory_wb_data_i[20] localMemory_wb_data_i[21]
+ localMemory_wb_data_i[22] localMemory_wb_data_i[23] localMemory_wb_data_i[24] localMemory_wb_data_i[25]
+ localMemory_wb_data_i[26] localMemory_wb_data_i[27] localMemory_wb_data_i[28] localMemory_wb_data_i[29]
+ localMemory_wb_data_i[2] localMemory_wb_data_i[30] localMemory_wb_data_i[31] localMemory_wb_data_i[3]
+ localMemory_wb_data_i[4] localMemory_wb_data_i[5] localMemory_wb_data_i[6] localMemory_wb_data_i[7]
+ localMemory_wb_data_i[8] localMemory_wb_data_i[9] localMemory_wb_data_o[0] localMemory_wb_data_o[10]
+ localMemory_wb_data_o[11] localMemory_wb_data_o[12] localMemory_wb_data_o[13] localMemory_wb_data_o[14]
+ localMemory_wb_data_o[15] localMemory_wb_data_o[16] localMemory_wb_data_o[17] localMemory_wb_data_o[18]
+ localMemory_wb_data_o[19] localMemory_wb_data_o[1] localMemory_wb_data_o[20] localMemory_wb_data_o[21]
+ localMemory_wb_data_o[22] localMemory_wb_data_o[23] localMemory_wb_data_o[24] localMemory_wb_data_o[25]
+ localMemory_wb_data_o[26] localMemory_wb_data_o[27] localMemory_wb_data_o[28] localMemory_wb_data_o[29]
+ localMemory_wb_data_o[2] localMemory_wb_data_o[30] localMemory_wb_data_o[31] localMemory_wb_data_o[3]
+ localMemory_wb_data_o[4] localMemory_wb_data_o[5] localMemory_wb_data_o[6] localMemory_wb_data_o[7]
+ localMemory_wb_data_o[8] localMemory_wb_data_o[9] localMemory_wb_error_o localMemory_wb_sel_i[0]
+ localMemory_wb_sel_i[1] localMemory_wb_sel_i[2] localMemory_wb_sel_i[3] localMemory_wb_stall_o
+ localMemory_wb_stb_i localMemory_wb_we_i manufacturerID[0] manufacturerID[10] manufacturerID[1]
+ manufacturerID[2] manufacturerID[3] manufacturerID[4] manufacturerID[5] manufacturerID[6]
+ manufacturerID[7] manufacturerID[8] manufacturerID[9] partID[0] partID[10] partID[11]
+ partID[12] partID[13] partID[14] partID[15] partID[1] partID[2] partID[3] partID[4]
+ partID[5] partID[6] partID[7] partID[8] partID[9] probe_env[0] probe_env[1] probe_jtagInstruction[0]
+ probe_jtagInstruction[1] probe_jtagInstruction[2] probe_jtagInstruction[3] probe_jtagInstruction[4]
+ probe_programCounter[0] probe_programCounter[10] probe_programCounter[11] probe_programCounter[12]
+ probe_programCounter[13] probe_programCounter[14] probe_programCounter[15] probe_programCounter[16]
+ probe_programCounter[17] probe_programCounter[18] probe_programCounter[19] probe_programCounter[1]
+ probe_programCounter[20] probe_programCounter[21] probe_programCounter[22] probe_programCounter[23]
+ probe_programCounter[24] probe_programCounter[25] probe_programCounter[26] probe_programCounter[27]
+ probe_programCounter[28] probe_programCounter[29] probe_programCounter[2] probe_programCounter[30]
+ probe_programCounter[31] probe_programCounter[3] probe_programCounter[4] probe_programCounter[5]
+ probe_programCounter[6] probe_programCounter[7] probe_programCounter[8] probe_programCounter[9]
+ probe_state vccd1 versionID[0] versionID[1] versionID[2] versionID[3] vssd1 wb_clk_i
+ wb_rst_i web0 wmask0[0] wmask0[1] wmask0[2] wmask0[3]
XFILLER_228_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09671_ _19039_/Q _19007_/Q _09671_/S vssd1 vssd1 vccd1 vccd1 _09671_/X sky130_fd_sc_hd__mux2_1
XFILLER_255_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18869_ _19055_/CLK _18869_/D vssd1 vssd1 vccd1 vccd1 _18869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ _09105_/A _11452_/A vssd1 vssd1 vccd1 vccd1 _09105_/X sky130_fd_sc_hd__or2_1
XFILLER_176_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09036_ _11691_/B1 _12409_/A2 _09035_/X _11692_/A1 _18392_/Q vssd1 vssd1 vccd1 vccd1
+ _09036_/X sky130_fd_sc_hd__o32a_1
XFILLER_191_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1807 _14442_/B vssd1 vssd1 vccd1 vccd1 _14451_/B sky130_fd_sc_hd__clkbuf_4
Xfanout820 _14307_/Y vssd1 vssd1 vccd1 vccd1 _14325_/S sky130_fd_sc_hd__buf_12
Xfanout1818 _17366_/A vssd1 vssd1 vccd1 vccd1 _17592_/B sky130_fd_sc_hd__buf_4
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout831 _16542_/A0 vssd1 vssd1 vccd1 vccd1 _16608_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout1829 _17326_/A vssd1 vssd1 vccd1 vccd1 _17419_/C1 sky130_fd_sc_hd__buf_4
X_09938_ _09936_/X _09937_/X _10265_/A vssd1 vssd1 vccd1 vccd1 _09938_/X sky130_fd_sc_hd__mux2_1
Xfanout842 _17678_/A0 vssd1 vssd1 vccd1 vccd1 _16611_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_89_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout853 _10792_/A2 vssd1 vssd1 vccd1 vccd1 _16547_/A0 sky130_fd_sc_hd__clkbuf_2
Xfanout864 _10341_/A2 vssd1 vssd1 vccd1 vccd1 _16619_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout875 _17721_/A0 vssd1 vssd1 vccd1 vccd1 _16522_/A0 sky130_fd_sc_hd__clkbuf_2
Xfanout886 _12943_/S vssd1 vssd1 vccd1 vccd1 _12933_/A sky130_fd_sc_hd__buf_6
Xfanout897 _09334_/X vssd1 vssd1 vccd1 vccd1 _16203_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09869_ _08901_/A _18135_/Q _18781_/Q _09885_/S _10747_/A1 vssd1 vssd1 vccd1 vccd1
+ _09869_/X sky130_fd_sc_hd__a221o_1
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _10121_/B _11845_/B _11952_/A2 vssd1 vssd1 vccd1 vccd1 _11903_/A sky130_fd_sc_hd__o21a_2
XFILLER_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12880_ _13039_/S _12877_/Y _12879_/Y _13354_/A vssd1 vssd1 vccd1 vccd1 _12880_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_202 _14164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _17906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11831_ _11844_/A _11831_/B vssd1 vssd1 vccd1 vccd1 _11831_/X sky130_fd_sc_hd__and2_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_224 _18383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _18393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 _18725_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_257 input205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 input227/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14576_/A _14550_/B vssd1 vssd1 vccd1 vccd1 _18383_/D sky130_fd_sc_hd__or2_1
XFILLER_214_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _18580_/Q _14349_/B _11769_/B1 _13545_/B vssd1 vssd1 vccd1 vccd1 _11762_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_279 input243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13501_ _19345_/Q _13950_/A2 _13950_/B1 _19473_/Q _13950_/C1 vssd1 vssd1 vccd1 vccd1
+ _13501_/X sky130_fd_sc_hd__a221o_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _09611_/A _10713_/A2 _11023_/B1 vssd1 vssd1 vccd1 vccd1 _10713_/X sky130_fd_sc_hd__o21a_1
X_14481_ _18333_/Q _17685_/A0 _14485_/S vssd1 vssd1 vccd1 vccd1 _18333_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11693_ _18203_/Q _11695_/B vssd1 vssd1 vccd1 vccd1 _11693_/Y sky130_fd_sc_hd__nand2_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16220_ _17717_/A0 _18836_/Q _16226_/S vssd1 vssd1 vccd1 vccd1 _18836_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13432_ _19343_/Q _13950_/A2 _13950_/B1 _19471_/Q _13950_/C1 vssd1 vssd1 vccd1 vccd1
+ _13432_/X sky130_fd_sc_hd__a221o_1
X_10644_ _10662_/A1 _19577_/Q _10645_/S _19609_/Q _10668_/S vssd1 vssd1 vccd1 vccd1
+ _10644_/X sky130_fd_sc_hd__o221a_1
XFILLER_139_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16151_ _16154_/A _16154_/B _16150_/X _16149_/A vssd1 vssd1 vccd1 vccd1 _16151_/X
+ sky130_fd_sc_hd__a31o_1
X_10575_ _19091_/Q _18995_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _10575_/X sky130_fd_sc_hd__mux2_1
X_13363_ _13363_/A vssd1 vssd1 vccd1 vccd1 _13363_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15102_ _17591_/A _17591_/B vssd1 vssd1 vccd1 vccd1 _15102_/Y sky130_fd_sc_hd__nor2_4
XFILLER_6_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12314_ _12315_/B _12314_/B vssd1 vssd1 vccd1 vccd1 _12314_/X sky130_fd_sc_hd__or2_4
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16082_ _16096_/A1 _16081_/Y _17725_/C1 vssd1 vssd1 vccd1 vccd1 _18743_/D sky130_fd_sc_hd__a21oi_1
XFILLER_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13294_ _13294_/A _13330_/B vssd1 vssd1 vccd1 vccd1 _13294_/X sky130_fd_sc_hd__or2_1
XFILLER_138_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15033_ _18522_/Q input199/X _15038_/S vssd1 vssd1 vccd1 vccd1 _18522_/D sky130_fd_sc_hd__mux2_1
X_12245_ _17881_/Q _12248_/C _12243_/A vssd1 vssd1 vccd1 vccd1 _12245_/Y sky130_fd_sc_hd__a21oi_1
X_12176_ _17855_/Q _17854_/Q _12176_/C vssd1 vssd1 vccd1 vccd1 _12178_/B sky130_fd_sc_hd__and3_1
XFILLER_122_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ _11125_/X _11126_/X _11127_/S vssd1 vssd1 vccd1 vccd1 _11127_/X sky130_fd_sc_hd__mux2_1
X_16984_ _17117_/B _17044_/A2 _16983_/X _17378_/A vssd1 vssd1 vccd1 vccd1 _19328_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15935_ input4/X input270/X _15947_/S vssd1 vssd1 vccd1 vccd1 _15935_/X sky130_fd_sc_hd__mux2_1
X_18723_ _18775_/CLK _18723_/D vssd1 vssd1 vccd1 vccd1 _18723_/Q sky130_fd_sc_hd__dfxtp_1
X_11058_ _11061_/B vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__inv_2
XFILLER_95_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19596_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10009_ _10009_/A _10009_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10009_/X sky130_fd_sc_hd__or3_2
X_18654_ _19624_/CLK _18654_/D vssd1 vssd1 vccd1 vccd1 _18654_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15866_ _15866_/A _15941_/S _15905_/C vssd1 vssd1 vccd1 vccd1 _15866_/X sky130_fd_sc_hd__and3_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14817_ _14813_/Y _14816_/X _14950_/B1 vssd1 vssd1 vccd1 vccd1 _14817_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17605_ _19382_/Q _15086_/B input183/X _17592_/X _17623_/B1 vssd1 vssd1 vccd1 vccd1
+ _17605_/X sky130_fd_sc_hd__a41o_1
XFILLER_92_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18585_ _19484_/CLK _18585_/D vssd1 vssd1 vccd1 vccd1 _18585_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_252_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ _15781_/S _15796_/Y _19487_/Q vssd1 vssd1 vccd1 vccd1 _15797_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17536_ _19518_/Q _17493_/B _17535_/X _17356_/A vssd1 vssd1 vccd1 vccd1 _19518_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_251_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14748_ _14745_/Y _14747_/Y _14879_/B1 vssd1 vssd1 vccd1 vccd1 _14748_/Y sky130_fd_sc_hd__a21oi_4
X_17467_ _18116_/Q _17545_/C1 _17465_/X _17466_/X vssd1 vssd1 vccd1 vccd1 _17467_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14679_ _14681_/C _14679_/B _14681_/B _14679_/D vssd1 vssd1 vccd1 vccd1 _14679_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19206_ _19206_/CLK _19206_/D vssd1 vssd1 vccd1 vccd1 _19206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16418_ _16418_/A0 _19027_/Q _16420_/S vssd1 vssd1 vccd1 vccd1 _19027_/D sky130_fd_sc_hd__mux2_1
X_17398_ _18102_/Q _17426_/B1 _17397_/X vssd1 vssd1 vccd1 vccd1 _17398_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_186_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19137_ _19147_/CLK _19137_/D vssd1 vssd1 vccd1 vccd1 _19137_/Q sky130_fd_sc_hd__dfxtp_1
X_16349_ _18961_/Q _16548_/A0 _16352_/S vssd1 vssd1 vccd1 vccd1 _18961_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19068_ _19587_/CLK _19068_/D vssd1 vssd1 vccd1 vccd1 _19068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput401 _11923_/X vssd1 vssd1 vccd1 vccd1 din0[3] sky130_fd_sc_hd__buf_4
Xoutput412 _18482_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[11] sky130_fd_sc_hd__buf_4
X_18019_ _19589_/CLK _18019_/D vssd1 vssd1 vccd1 vccd1 _18019_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput423 _18492_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[21] sky130_fd_sc_hd__buf_4
XFILLER_161_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput434 _18502_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[31] sky130_fd_sc_hd__buf_4
Xoutput445 _18733_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[0] sky130_fd_sc_hd__buf_4
Xoutput456 _18116_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[15] sky130_fd_sc_hd__buf_4
Xoutput467 _18126_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[25] sky130_fd_sc_hd__buf_4
XFILLER_271_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput478 _18107_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[6] sky130_fd_sc_hd__buf_4
XFILLER_114_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09723_ _09721_/X _09722_/X _09723_/S vssd1 vssd1 vccd1 vccd1 _09723_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09654_ _18385_/Q _09656_/B1 _09331_/A _09653_/Y vssd1 vssd1 vccd1 vccd1 _09660_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_243_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ _10373_/S _09585_/B vssd1 vssd1 vccd1 vccd1 _09585_/X sky130_fd_sc_hd__or2_1
XFILLER_103_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10360_ _10366_/A1 _19222_/Q _19190_/Q _10370_/S _12766_/A0 vssd1 vssd1 vccd1 vccd1
+ _10360_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ _09245_/A _09028_/B vssd1 vssd1 vccd1 vccd1 _09019_/Y sky130_fd_sc_hd__nor2_2
X_10291_ _10289_/X _10290_/X _10300_/S vssd1 vssd1 vccd1 vccd1 _10291_/X sky130_fd_sc_hd__mux2_1
XFILLER_275_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12030_ _17890_/Q _12035_/B _12029_/Y _12383_/C1 vssd1 vssd1 vccd1 vccd1 _17792_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1604 _15104_/X vssd1 vssd1 vccd1 vccd1 _17550_/A sky130_fd_sc_hd__buf_4
XFILLER_120_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1615 _11707_/X vssd1 vssd1 vccd1 vccd1 _11711_/A sky130_fd_sc_hd__buf_6
Xfanout1626 _09908_/B1 vssd1 vssd1 vccd1 vccd1 _09656_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1637 _08858_/Y vssd1 vssd1 vccd1 vccd1 _12420_/A1 sky130_fd_sc_hd__buf_8
Xfanout650 _17045_/B vssd1 vssd1 vccd1 vccd1 _17041_/B sky130_fd_sc_hd__buf_4
Xfanout1648 _11618_/A1 vssd1 vssd1 vccd1 vccd1 _11277_/A1 sky130_fd_sc_hd__buf_6
Xfanout1659 _11506_/A1 vssd1 vssd1 vccd1 vccd1 _11513_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout661 _13781_/A2 vssd1 vssd1 vccd1 vccd1 _13947_/A2 sky130_fd_sc_hd__buf_4
Xfanout672 _14875_/A1 vssd1 vssd1 vccd1 vccd1 _14865_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_59_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13981_ _17955_/Q _14004_/A _13980_/Y _13981_/C1 vssd1 vssd1 vccd1 vccd1 _17955_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout683 _12570_/C vssd1 vssd1 vccd1 vccd1 _13950_/C1 sky130_fd_sc_hd__buf_6
Xfanout694 _13950_/A2 vssd1 vssd1 vccd1 vccd1 _13883_/A2 sky130_fd_sc_hd__buf_6
XFILLER_246_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15720_ _18129_/Q _15763_/A2 _15719_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _15722_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ _13314_/S _12932_/B vssd1 vssd1 vccd1 vccd1 _12932_/X sky130_fd_sc_hd__or2_1
XFILLER_58_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15651_ _15651_/A _15651_/B vssd1 vssd1 vccd1 vccd1 _15653_/A sky130_fd_sc_hd__nand2_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _17825_/Q _12862_/X _13944_/B vssd1 vssd1 vccd1 vccd1 _12863_/X sky130_fd_sc_hd__mux2_2
XFILLER_206_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _17694_/A0 _18409_/Q _14622_/S vssd1 vssd1 vccd1 vccd1 _18409_/D sky130_fd_sc_hd__mux2_1
X_18370_ _19648_/CLK _18370_/D vssd1 vssd1 vccd1 vccd1 _18370_/Q sky130_fd_sc_hd__dfxtp_1
X_11814_ _11818_/A _11818_/B _11814_/C vssd1 vssd1 vccd1 vccd1 _11814_/X sky130_fd_sc_hd__and3_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15582_ _18582_/Q _15581_/C _18583_/Q vssd1 vssd1 vccd1 vccd1 _15583_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12693_/X _12697_/X _12818_/S vssd1 vssd1 vccd1 vccd1 _12794_/X sky130_fd_sc_hd__mux2_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _19458_/Q _17563_/A _17377_/S vssd1 vssd1 vccd1 vccd1 _17322_/B sky130_fd_sc_hd__mux2_1
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _18375_/Q _14559_/A2 _14559_/B1 input32/X vssd1 vssd1 vccd1 vccd1 _14534_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _13127_/A sky130_fd_sc_hd__nor2_8
XFILLER_144_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17252_ _17250_/Y _17251_/X _17338_/A vssd1 vssd1 vccd1 vccd1 _19434_/D sky130_fd_sc_hd__o21a_1
X_14464_ _18316_/Q _17701_/A0 _14485_/S vssd1 vssd1 vccd1 vccd1 _18316_/D sky130_fd_sc_hd__mux2_1
X_11676_ _11676_/A _11676_/B vssd1 vssd1 vccd1 vccd1 _13512_/B sky130_fd_sc_hd__xnor2_4
X_16203_ _16203_/A0 _18819_/Q _16222_/S vssd1 vssd1 vccd1 vccd1 _18819_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13415_ _13135_/S _13131_/X _13136_/S vssd1 vssd1 vccd1 vccd1 _13415_/Y sky130_fd_sc_hd__a21oi_1
X_17183_ _17210_/A _17183_/B vssd1 vssd1 vccd1 vccd1 _19412_/D sky130_fd_sc_hd__nor2_1
X_10627_ _10625_/X _10626_/X _10632_/S vssd1 vssd1 vccd1 vccd1 _10627_/X sky130_fd_sc_hd__mux2_1
X_14395_ _16470_/A0 _18246_/Q _14415_/S vssd1 vssd1 vccd1 vccd1 _18246_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16134_ _16142_/A1 _16133_/Y _16142_/B1 vssd1 vssd1 vccd1 vccd1 _18769_/D sky130_fd_sc_hd__a21oi_1
X_13346_ _13637_/A _14000_/B _13333_/Y vssd1 vssd1 vccd1 vccd1 _13346_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10558_ _10633_/A _10558_/B vssd1 vssd1 vccd1 vccd1 _10558_/X sky130_fd_sc_hd__or2_1
XFILLER_255_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16065_ _16056_/Y _16075_/B _16063_/Y _16064_/X vssd1 vssd1 vccd1 vccd1 _16065_/Y
+ sky130_fd_sc_hd__a31oi_1
X_13277_ _19533_/Q _19501_/Q _13277_/S vssd1 vssd1 vccd1 vccd1 _13277_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10489_ _11103_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10489_/Y sky130_fd_sc_hd__nor2_1
X_15016_ _18505_/Q input201/X _16627_/S vssd1 vssd1 vccd1 vccd1 _18505_/D sky130_fd_sc_hd__mux2_1
X_12228_ _17874_/Q _12226_/B _12227_/Y vssd1 vssd1 vccd1 vccd1 _17874_/D sky130_fd_sc_hd__o21a_1
XFILLER_151_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12159_ _17848_/Q _12160_/C _17849_/Q vssd1 vssd1 vccd1 vccd1 _12161_/B sky130_fd_sc_hd__a21oi_1
XFILLER_284_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16967_ _19326_/Q _17211_/B _16967_/S vssd1 vssd1 vccd1 vccd1 _16968_/B sky130_fd_sc_hd__mux2_1
XFILLER_272_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18706_ _19306_/CLK _18706_/D vssd1 vssd1 vccd1 vccd1 _18706_/Q sky130_fd_sc_hd__dfxtp_1
X_15918_ _18681_/Q _15918_/A2 _15948_/C1 _15917_/X vssd1 vssd1 vccd1 vccd1 _15918_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_265_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16898_ _16898_/A1 _17933_/Q _16897_/X vssd1 vssd1 vccd1 vccd1 _17585_/A sky130_fd_sc_hd__o21a_4
XFILLER_64_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18637_ _19076_/CLK _18637_/D vssd1 vssd1 vccd1 vccd1 _18637_/Q sky130_fd_sc_hd__dfxtp_4
X_15849_ _15849_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15955_/B sky130_fd_sc_hd__or2_4
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09370_ _18851_/Q _18883_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09370_/X sky130_fd_sc_hd__mux2_1
X_18568_ _19525_/CLK _18568_/D vssd1 vssd1 vccd1 vccd1 _18568_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_252_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17519_ _19515_/Q _17517_/B _17518_/X _17368_/A vssd1 vssd1 vccd1 vccd1 _19515_/D
+ sky130_fd_sc_hd__o211a_1
X_18499_ _18501_/CLK _18499_/D vssd1 vssd1 vccd1 vccd1 _18499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput286 _11961_/X vssd1 vssd1 vccd1 vccd1 addr0[1] sky130_fd_sc_hd__buf_4
Xoutput297 _11913_/X vssd1 vssd1 vccd1 vccd1 addr1[3] sky130_fd_sc_hd__buf_4
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09706_ _09702_/X _09703_/X _10300_/S vssd1 vssd1 vccd1 vccd1 _09706_/X sky130_fd_sc_hd__mux2_1
XFILLER_244_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09637_ _19623_/Q _18912_/Q _10687_/S vssd1 vssd1 vccd1 vccd1 _09637_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ _18386_/Q _09656_/B1 _09331_/A _09567_/Y vssd1 vssd1 vccd1 vccd1 _09574_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09499_ _09497_/X _09498_/X _09723_/S vssd1 vssd1 vccd1 vccd1 _09499_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11530_ _11215_/B _11677_/B _13468_/S vssd1 vssd1 vccd1 vccd1 _11676_/B sky130_fd_sc_hd__o21bai_4
XFILLER_211_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11461_ _18419_/Q _11479_/B _11460_/X _10403_/S vssd1 vssd1 vccd1 vccd1 _11461_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13200_ _18110_/Q _13201_/B vssd1 vssd1 vccd1 vccd1 _13271_/C sky130_fd_sc_hd__and2_2
X_10412_ _10409_/X _10411_/X _10405_/X vssd1 vssd1 vccd1 vccd1 _10412_/Y sky130_fd_sc_hd__a21oi_4
X_11392_ _19631_/Q _18920_/Q _11477_/S vssd1 vssd1 vccd1 vccd1 _11392_/X sky130_fd_sc_hd__mux2_1
X_14180_ _18701_/Q _18088_/Q _14186_/S vssd1 vssd1 vccd1 vccd1 _14181_/B sky130_fd_sc_hd__mux2_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _13130_/A _12934_/Y _13130_/Y vssd1 vssd1 vccd1 vccd1 _13131_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10343_ _17915_/Q _11441_/B _11489_/B1 _10342_/Y vssd1 vssd1 vccd1 vccd1 _10381_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_180_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10274_ _18560_/Q _18435_/Q _10299_/S vssd1 vssd1 vccd1 vccd1 _10274_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13062_ _08818_/Y _13246_/B1 _12570_/C vssd1 vssd1 vccd1 vccd1 _13062_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12013_ _17780_/Q _16548_/A0 _12013_/S vssd1 vssd1 vccd1 vccd1 _17780_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17870_ _19310_/CLK _17870_/D vssd1 vssd1 vccd1 vccd1 _17870_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1401 _09542_/S vssd1 vssd1 vccd1 vccd1 _11160_/S sky130_fd_sc_hd__buf_6
Xfanout1412 fanout1415/X vssd1 vssd1 vccd1 vccd1 _09179_/B sky130_fd_sc_hd__buf_6
Xfanout1423 _11379_/S vssd1 vssd1 vccd1 vccd1 _11462_/S sky130_fd_sc_hd__buf_4
XFILLER_215_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1434 _10557_/S vssd1 vssd1 vccd1 vccd1 _10784_/S sky130_fd_sc_hd__buf_6
XFILLER_120_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1445 _11002_/C1 vssd1 vssd1 vccd1 vccd1 _10408_/S sky130_fd_sc_hd__buf_4
X_16821_ _16821_/A _17813_/Q vssd1 vssd1 vccd1 vccd1 _16840_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1456 _10337_/S1 vssd1 vssd1 vccd1 vccd1 _09136_/S sky130_fd_sc_hd__buf_4
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1467 fanout1469/X vssd1 vssd1 vccd1 vccd1 _11604_/S sky130_fd_sc_hd__buf_6
Xfanout1478 _09801_/S vssd1 vssd1 vccd1 vccd1 _11613_/S sky130_fd_sc_hd__buf_6
XFILLER_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout491 _14889_/B1 vssd1 vssd1 vccd1 vccd1 _14720_/A sky130_fd_sc_hd__buf_4
Xfanout1489 fanout1525/X vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__clkbuf_4
X_16752_ _16752_/A _16752_/B _16754_/B vssd1 vssd1 vccd1 vccd1 _19270_/D sky130_fd_sc_hd__nor3_1
X_19540_ _19540_/CLK _19540_/D vssd1 vssd1 vccd1 vccd1 _19540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13964_ _11628_/A _13962_/Y _13963_/Y vssd1 vssd1 vccd1 vccd1 _13964_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_234_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15703_ _15689_/A _15689_/B _15684_/B vssd1 vssd1 vccd1 vccd1 _15707_/B sky130_fd_sc_hd__a21oi_1
X_12915_ _12580_/A _12576_/B _12584_/Y input4/X vssd1 vssd1 vccd1 vccd1 _12915_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_262_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16683_ _19240_/Q _19237_/Q _16683_/C _16683_/D vssd1 vssd1 vccd1 vccd1 _16690_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19471_ _19471_/CLK _19471_/D vssd1 vssd1 vccd1 vccd1 _19471_/Q sky130_fd_sc_hd__dfxtp_1
X_13895_ _13891_/A _12837_/B _13962_/B _11634_/A _13894_/Y vssd1 vssd1 vccd1 vccd1
+ _13895_/X sky130_fd_sc_hd__o221a_1
XFILLER_250_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15634_ _18585_/Q _15718_/A2 _15633_/X _17374_/A vssd1 vssd1 vccd1 vccd1 _18585_/D
+ sky130_fd_sc_hd__o211a_1
X_18422_ _19601_/CLK _18422_/D vssd1 vssd1 vccd1 vccd1 _18422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ _13100_/A _12846_/B vssd1 vssd1 vccd1 vccd1 _17921_/D sky130_fd_sc_hd__and2_1
XFILLER_261_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _19631_/CLK _18353_/D vssd1 vssd1 vccd1 vccd1 _18353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15565_ _15560_/X _15563_/X _15564_/Y vssd1 vssd1 vccd1 vccd1 _15565_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12777_ _19297_/Q _12583_/Y _12584_/Y input2/X _12776_/X vssd1 vssd1 vccd1 vccd1
+ _12777_/X sky130_fd_sc_hd__a221o_4
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17304_ _19452_/Q _17307_/B vssd1 vssd1 vccd1 vccd1 _17304_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14516_ _16618_/A0 _18366_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _18366_/D sky130_fd_sc_hd__mux2_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11728_ _11728_/A _13904_/B _11728_/C vssd1 vssd1 vccd1 vccd1 _15039_/B sky130_fd_sc_hd__and3_4
X_18284_ _18778_/CLK _18284_/D vssd1 vssd1 vccd1 vccd1 _18284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15496_ _15496_/A _15496_/B vssd1 vssd1 vccd1 vccd1 _15497_/B sky130_fd_sc_hd__nand2_1
XFILLER_230_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17235_ _19429_/Q _17256_/B vssd1 vssd1 vccd1 vccd1 _17235_/Y sky130_fd_sc_hd__nand2_1
X_14447_ _18586_/Q _14450_/B vssd1 vssd1 vccd1 vccd1 _18299_/D sky130_fd_sc_hd__and2_1
XFILLER_175_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11659_ _12740_/B _11832_/B _14141_/A vssd1 vssd1 vccd1 vccd1 _11659_/X sky130_fd_sc_hd__mux2_1
XFILLER_266_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17166_ _17166_/A _17589_/A vssd1 vssd1 vccd1 vccd1 _17468_/A sky130_fd_sc_hd__nand2_1
X_14378_ _18230_/Q _17685_/A0 _14382_/S vssd1 vssd1 vccd1 vccd1 _18230_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16117_ _18761_/Q _16139_/B vssd1 vssd1 vccd1 vccd1 _16117_/Y sky130_fd_sc_hd__nand2_1
XFILLER_171_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13329_ _13937_/A _13329_/B vssd1 vssd1 vccd1 vccd1 _13329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17097_ _19382_/Q _17107_/B vssd1 vssd1 vccd1 vccd1 _17097_/X sky130_fd_sc_hd__or2_1
XFILLER_171_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16048_ _16048_/A _16048_/B vssd1 vssd1 vccd1 vccd1 _18735_/D sky130_fd_sc_hd__or2_1
XFILLER_115_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08870_ _08870_/A _12443_/A _12438_/B vssd1 vssd1 vccd1 vccd1 _12435_/A sky130_fd_sc_hd__or3_4
XFILLER_97_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17999_ _19601_/CLK _17999_/D vssd1 vssd1 vccd1 vccd1 _17999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09422_ _09420_/X _09421_/X _09429_/S vssd1 vssd1 vccd1 vccd1 _09422_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09353_ _18634_/Q _11395_/C vssd1 vssd1 vccd1 vccd1 _09353_/X sky130_fd_sc_hd__or2_1
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09284_ _12389_/A1 _09282_/X _09283_/X _12962_/A0 vssd1 vssd1 vccd1 vccd1 _09284_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_193_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08999_ _08999_/A _11218_/A vssd1 vssd1 vccd1 vccd1 _10309_/A sky130_fd_sc_hd__nor2_1
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_188_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19155_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_229_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_117_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19261_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_216_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10961_ _10959_/X _10960_/X _11127_/S vssd1 vssd1 vccd1 vccd1 _10961_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12700_ _12692_/X _12699_/X _13039_/S vssd1 vssd1 vccd1 vccd1 _12700_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13680_ _17846_/Q _13744_/A2 _13744_/B1 _17878_/Q vssd1 vssd1 vccd1 vccd1 _13680_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10892_ _11358_/A _10891_/X _11608_/C1 vssd1 vssd1 vccd1 vccd1 _10892_/X sky130_fd_sc_hd__a21o_1
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12631_ _13465_/B _13465_/C _13465_/A vssd1 vssd1 vccd1 vccd1 _13466_/A sky130_fd_sc_hd__a21oi_4
XPHY_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15350_ _15340_/Y _15344_/Y _15349_/Y vssd1 vssd1 vccd1 vccd1 _15350_/Y sky130_fd_sc_hd__o21ai_1
XPHY_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12562_ _12580_/A _12562_/B vssd1 vssd1 vccd1 vccd1 _12562_/X sky130_fd_sc_hd__or2_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14301_ _16619_/A0 _18160_/Q _14301_/S vssd1 vssd1 vccd1 vccd1 _18160_/D sky130_fd_sc_hd__mux2_1
X_11513_ _11513_/A1 _18606_/Q _18177_/Q _11513_/B2 vssd1 vssd1 vccd1 vccd1 _11513_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15281_ _19464_/Q _15280_/X _15400_/S vssd1 vssd1 vccd1 vccd1 _15281_/X sky130_fd_sc_hd__mux2_1
X_12493_ _12488_/A _17915_/Q _12492_/X vssd1 vssd1 vccd1 vccd1 _12554_/B sky130_fd_sc_hd__a21o_4
XFILLER_200_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17020_ _17175_/B _17046_/A2 _17019_/X _17354_/A vssd1 vssd1 vccd1 vccd1 _19346_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14232_ _18114_/Q _14260_/B vssd1 vssd1 vccd1 vccd1 _14232_/X sky130_fd_sc_hd__or2_1
X_11444_ _12597_/A _11445_/B vssd1 vssd1 vccd1 vccd1 _13357_/S sky130_fd_sc_hd__and2_4
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14163_ _14164_/B _15953_/A vssd1 vssd1 vccd1 vccd1 _16143_/B sky130_fd_sc_hd__nor2_1
X_11375_ _17933_/Q _11451_/A2 _11374_/X _11451_/B2 vssd1 vssd1 vccd1 vccd1 _11375_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_153_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13114_ input261/X _12506_/X _13103_/X _13113_/X _12510_/X vssd1 vssd1 vccd1 vccd1
+ _13116_/A sky130_fd_sc_hd__o221a_1
X_10326_ _10326_/A _10326_/B vssd1 vssd1 vccd1 vccd1 _10326_/Y sky130_fd_sc_hd__nand2_1
X_14094_ _17677_/A0 _18034_/Q _14106_/S vssd1 vssd1 vccd1 vccd1 _18034_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18971_ _19195_/CLK _18971_/D vssd1 vssd1 vccd1 vccd1 _18971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13045_ _13358_/A1 _13044_/X _09648_/B vssd1 vssd1 vccd1 vccd1 _13045_/X sky130_fd_sc_hd__a21o_2
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17922_ _17930_/CLK _17922_/D vssd1 vssd1 vccd1 vccd1 _17922_/Q sky130_fd_sc_hd__dfxtp_4
X_10257_ _10263_/A1 _19582_/Q _10253_/C _19614_/Q vssd1 vssd1 vccd1 vccd1 _10257_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1220 _12762_/A vssd1 vssd1 vccd1 vccd1 _12448_/C sky130_fd_sc_hd__buf_8
XFILLER_121_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1231 _14692_/A2 vssd1 vssd1 vccd1 vccd1 _12305_/B1 sky130_fd_sc_hd__buf_6
XFILLER_67_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10188_ _10334_/A1 _19160_/Q _10090_/S _19128_/Q vssd1 vssd1 vccd1 vccd1 _10188_/X
+ sky130_fd_sc_hd__o22a_1
X_17853_ _19327_/CLK _17853_/D vssd1 vssd1 vccd1 vccd1 _17853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1242 _09042_/Y vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__buf_4
XFILLER_267_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1253 _10905_/S vssd1 vssd1 vccd1 vccd1 _11337_/B sky130_fd_sc_hd__buf_4
XFILLER_227_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1264 _08890_/Y vssd1 vssd1 vccd1 vccd1 _13938_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_266_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16804_ _19290_/Q _16807_/C _16812_/B1 vssd1 vssd1 vccd1 vccd1 _16804_/Y sky130_fd_sc_hd__o21ai_1
Xfanout1275 _12264_/X vssd1 vssd1 vccd1 vccd1 _13260_/A sky130_fd_sc_hd__buf_8
Xfanout1286 _15854_/B vssd1 vssd1 vccd1 vccd1 _15970_/A2 sky130_fd_sc_hd__buf_6
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17784_ _19612_/CLK _17784_/D vssd1 vssd1 vccd1 vccd1 _17784_/Q sky130_fd_sc_hd__dfxtp_1
X_14996_ _14996_/A1 _14995_/X _11715_/B vssd1 vssd1 vccd1 vccd1 _14996_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_66_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1297 _14586_/A vssd1 vssd1 vccd1 vccd1 _14576_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_254_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19523_ _19525_/CLK _19523_/D vssd1 vssd1 vccd1 vccd1 _19523_/Q sky130_fd_sc_hd__dfxtp_1
X_16735_ _16737_/A _16735_/B _16739_/C vssd1 vssd1 vccd1 vccd1 _19264_/D sky130_fd_sc_hd__nor3_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13947_ _19521_/Q _13947_/A2 _13947_/B1 _13946_/X vssd1 vssd1 vccd1 vccd1 _13947_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16666_ _19244_/Q _19243_/Q _19242_/Q _19241_/Q vssd1 vssd1 vccd1 vccd1 _16677_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_250_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19454_ _19507_/CLK _19454_/D vssd1 vssd1 vccd1 vccd1 _19454_/Q sky130_fd_sc_hd__dfxtp_4
X_13878_ _17884_/Q _13945_/A2 _13877_/X _13920_/B2 vssd1 vssd1 vccd1 vccd1 _13878_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15617_ _14252_/A _15763_/A2 _15616_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _15618_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18405_ _19477_/CLK _18405_/D vssd1 vssd1 vccd1 vccd1 _18405_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12829_ _12808_/X _12828_/X _13136_/S vssd1 vssd1 vccd1 vccd1 _13911_/B sky130_fd_sc_hd__mux2_4
X_16597_ _16597_/A0 _19200_/Q _16619_/S vssd1 vssd1 vccd1 vccd1 _19200_/D sky130_fd_sc_hd__mux2_1
X_19385_ _19481_/CLK _19385_/D vssd1 vssd1 vccd1 vccd1 _19385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18336_ _19615_/CLK _18336_/D vssd1 vssd1 vccd1 vccd1 _18336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15548_ _15549_/A _15623_/A vssd1 vssd1 vccd1 vccd1 _15764_/A sky130_fd_sc_hd__and2_1
XFILLER_231_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18267_ _19639_/CLK _18267_/D vssd1 vssd1 vccd1 vccd1 _18267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15479_ _15502_/B _13482_/Y _15133_/B _15478_/Y vssd1 vssd1 vccd1 vccd1 _15479_/X
+ sky130_fd_sc_hd__a31o_1
X_17218_ _17250_/B vssd1 vssd1 vccd1 vccd1 _17219_/B sky130_fd_sc_hd__inv_2
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18198_ _18817_/CLK _18198_/D vssd1 vssd1 vccd1 vccd1 _18198_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17149_ _19401_/Q fanout534/X _17438_/A _17212_/B2 vssd1 vssd1 vccd1 vccd1 _17150_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09971_ _19100_/Q _19132_/Q _09973_/S vssd1 vssd1 vccd1 vccd1 _09971_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08922_ _12089_/A _17797_/Q vssd1 vssd1 vccd1 vccd1 _14074_/C sky130_fd_sc_hd__nand2_8
XFILLER_257_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08853_ _17896_/Q vssd1 vssd1 vccd1 vccd1 _08853_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09405_ _14220_/A _13185_/A vssd1 vssd1 vccd1 vccd1 _09405_/Y sky130_fd_sc_hd__nand2_2
XFILLER_213_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09336_ _18851_/Q _18883_/Q _09937_/S vssd1 vssd1 vccd1 vccd1 _09336_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09267_ _18635_/Q _09269_/S vssd1 vssd1 vccd1 vccd1 _09267_/X sky130_fd_sc_hd__or2_1
XFILLER_193_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09198_ _18604_/Q _18175_/Q _10141_/S vssd1 vssd1 vccd1 vccd1 _09198_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11160_ _19634_/Q _18923_/Q _11160_/S vssd1 vssd1 vccd1 vccd1 _11160_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10111_ _10250_/S _10106_/X _10110_/X vssd1 vssd1 vccd1 vccd1 _10111_/Y sky130_fd_sc_hd__o21ai_2
X_11091_ _18253_/Q _10929_/S _10785_/A _11090_/X vssd1 vssd1 vccd1 vccd1 _11091_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_283_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _10036_/S _10029_/X _10030_/X vssd1 vssd1 vccd1 vccd1 _10042_/Y sky130_fd_sc_hd__o21ai_1
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14850_ _14912_/A1 _13459_/Y _15003_/B1 _18642_/Q _15003_/C1 vssd1 vssd1 vccd1 vccd1
+ _14850_/X sky130_fd_sc_hd__a221o_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _12444_/X _13800_/Y _13792_/X vssd1 vssd1 vccd1 vccd1 _13801_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14781_ _14779_/X _14780_/X _14964_/B1 vssd1 vssd1 vccd1 vccd1 _14781_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11993_ _17760_/Q _17694_/A0 _12013_/S vssd1 vssd1 vccd1 vccd1 _17760_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16520_ _16553_/A0 _19126_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _19126_/D sky130_fd_sc_hd__mux2_1
XFILLER_217_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13732_ _12732_/S _13137_/Y _13140_/X _13896_/B2 vssd1 vssd1 vccd1 vccd1 _13732_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10944_ _10917_/X _10920_/X _10399_/A vssd1 vssd1 vccd1 vccd1 _10944_/X sky130_fd_sc_hd__a21o_1
XFILLER_205_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16451_ _19059_/Q _17716_/A0 _16453_/S vssd1 vssd1 vccd1 vccd1 _19059_/D sky130_fd_sc_hd__mux2_1
X_13663_ _13676_/B _13761_/B vssd1 vssd1 vccd1 vccd1 _13663_/X sky130_fd_sc_hd__or2_1
XFILLER_232_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10875_ _18256_/Q _18831_/Q _18459_/Q _18360_/Q _11604_/S _11357_/S1 vssd1 vssd1
+ vccd1 vccd1 _10876_/B sky130_fd_sc_hd__mux4_1
XFILLER_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15402_ _18575_/Q _15447_/B _15394_/X _15401_/X _17469_/C1 vssd1 vssd1 vccd1 vccd1
+ _18575_/D sky130_fd_sc_hd__o221a_1
X_19170_ _19625_/CLK _19170_/D vssd1 vssd1 vccd1 vccd1 _19170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _09647_/B _12614_/B vssd1 vssd1 vccd1 vccd1 _13083_/B sky130_fd_sc_hd__nand2b_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _16548_/A0 _18993_/Q _16385_/S vssd1 vssd1 vccd1 vccd1 _18993_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13594_ _14014_/B vssd1 vssd1 vccd1 vccd1 _13594_/Y sky130_fd_sc_hd__inv_2
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17901_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18121_ _18593_/CLK _18121_/D vssd1 vssd1 vccd1 vccd1 _18121_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ _15404_/B _13273_/Y _15381_/A3 _15332_/X vssd1 vssd1 vccd1 vccd1 _15333_/X
+ sky130_fd_sc_hd__a31o_1
X_12545_ _12545_/A _12579_/A vssd1 vssd1 vccd1 vccd1 _12545_/Y sky130_fd_sc_hd__nor2_4
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19146_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18052_ _19592_/CLK _18052_/D vssd1 vssd1 vccd1 vccd1 _18052_/Q sky130_fd_sc_hd__dfxtp_1
X_15264_ _08840_/Y _15307_/B _15243_/A _15242_/X _15218_/Y vssd1 vssd1 vccd1 vccd1
+ _15264_/Y sky130_fd_sc_hd__o32ai_4
X_12476_ _12483_/A _12476_/B vssd1 vssd1 vccd1 vccd1 _12476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17003_ _19338_/Q _17003_/B vssd1 vssd1 vccd1 vccd1 _17003_/X sky130_fd_sc_hd__or2_1
X_14215_ _18279_/Q _14252_/B _14214_/X _16046_/A vssd1 vssd1 vccd1 vccd1 _18105_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11427_ _11425_/X _11426_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _11428_/B sky130_fd_sc_hd__mux2_1
XANTENNA_5 _18200_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _15259_/B _13030_/Y _15285_/A3 _15194_/Y vssd1 vssd1 vccd1 vccd1 _15195_/X
+ sky130_fd_sc_hd__a31o_1
X_14146_ _14146_/A _14146_/B _14146_/C vssd1 vssd1 vccd1 vccd1 _14147_/D sky130_fd_sc_hd__or3_1
X_11358_ _11358_/A _11358_/B vssd1 vssd1 vccd1 vccd1 _11358_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10309_ _10309_/A _10309_/B vssd1 vssd1 vccd1 vccd1 _10309_/Y sky130_fd_sc_hd__nor2_1
X_14077_ _16593_/A0 _18017_/Q _14104_/S vssd1 vssd1 vccd1 vccd1 _18017_/D sky130_fd_sc_hd__mux2_1
X_18954_ _19146_/CLK _18954_/D vssd1 vssd1 vccd1 vccd1 _18954_/Q sky130_fd_sc_hd__dfxtp_1
X_11289_ _11133_/B2 _11288_/X _17641_/A0 _11624_/A1 vssd1 vssd1 vccd1 vccd1 _15426_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_267_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17905_ _19595_/CLK _17905_/D vssd1 vssd1 vccd1 vccd1 _17905_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13028_ _18106_/Q _14214_/A _13028_/C vssd1 vssd1 vccd1 vccd1 _13055_/B sky130_fd_sc_hd__and3_1
XFILLER_39_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18885_ _19203_/CLK _18885_/D vssd1 vssd1 vccd1 vccd1 _18885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1050 _17528_/B vssd1 vssd1 vccd1 vccd1 _17463_/A2 sky130_fd_sc_hd__buf_2
XFILLER_227_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1061 _13483_/B vssd1 vssd1 vccd1 vccd1 _13349_/B sky130_fd_sc_hd__buf_4
X_17836_ _19310_/CLK _17836_/D vssd1 vssd1 vccd1 vccd1 _17836_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1072 _14027_/A2 vssd1 vssd1 vccd1 vccd1 _14028_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_120_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1083 _09980_/A2 vssd1 vssd1 vccd1 vccd1 _17660_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1094 _11624_/A1 vssd1 vssd1 vccd1 vccd1 _11365_/B2 sky130_fd_sc_hd__buf_6
XFILLER_187_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17767_ _19595_/CLK _17767_/D vssd1 vssd1 vccd1 vccd1 _17767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14979_ _14979_/A1 _18272_/Q _14978_/Y _11712_/A vssd1 vssd1 vccd1 vccd1 _14979_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_47_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19506_ _19506_/CLK _19506_/D vssd1 vssd1 vccd1 vccd1 _19506_/Q sky130_fd_sc_hd__dfxtp_1
X_16718_ _19258_/Q _16715_/B _16716_/Y vssd1 vssd1 vccd1 vccd1 _19258_/D sky130_fd_sc_hd__o21a_1
XFILLER_223_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17698_ _17698_/A0 _19624_/Q _17719_/S vssd1 vssd1 vccd1 vccd1 _19624_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19437_ _19537_/CLK _19437_/D vssd1 vssd1 vccd1 vccd1 _19437_/Q sky130_fd_sc_hd__dfxtp_1
X_16649_ _19239_/Q _19238_/Q _16649_/C vssd1 vssd1 vccd1 vccd1 _16658_/C sky130_fd_sc_hd__and3_1
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19368_ _19464_/CLK _19368_/D vssd1 vssd1 vccd1 vccd1 _19368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09121_ _18027_/Q _17995_/Q _11455_/S vssd1 vssd1 vccd1 vccd1 _09121_/X sky130_fd_sc_hd__mux2_1
X_18319_ _19612_/CLK _18319_/D vssd1 vssd1 vccd1 vccd1 _18319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19299_ _19326_/CLK _19299_/D vssd1 vssd1 vccd1 vccd1 _19299_/Q sky130_fd_sc_hd__dfxtp_1
X_09052_ _11687_/A _09052_/B vssd1 vssd1 vccd1 vccd1 _09052_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09954_ _18876_/Q _10364_/B vssd1 vssd1 vccd1 vccd1 _09954_/X sky130_fd_sc_hd__or2_1
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08905_ _08932_/A _12053_/A _12051_/A vssd1 vssd1 vccd1 vccd1 _08905_/X sky130_fd_sc_hd__or3b_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09885_ _19101_/Q _19133_/Q _09885_/S vssd1 vssd1 vccd1 vccd1 _09885_/X sky130_fd_sc_hd__mux2_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _12461_/A vssd1 vssd1 vccd1 vccd1 _12460_/A sky130_fd_sc_hd__inv_6
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_406 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_417 _11845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_428 _11836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_439 _13096_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ _10658_/X _10659_/X _10668_/S vssd1 vssd1 vccd1 vccd1 _10660_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09319_ _13188_/A vssd1 vssd1 vccd1 vccd1 _11750_/A sky130_fd_sc_hd__inv_2
XFILLER_22_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10591_ _18463_/Q _18364_/Q _10667_/S vssd1 vssd1 vccd1 vccd1 _10591_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12330_ _17817_/Q _17816_/Q _12330_/C _12330_/D vssd1 vssd1 vccd1 vccd1 _12333_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_194_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12261_ _17894_/Q _12261_/B vssd1 vssd1 vccd1 vccd1 _12315_/B sky130_fd_sc_hd__nand2_2
XFILLER_5_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14000_ _14032_/B _14000_/B vssd1 vssd1 vccd1 vccd1 _14000_/Y sky130_fd_sc_hd__nand2_1
X_11212_ _11214_/B vssd1 vssd1 vccd1 vccd1 _11212_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12192_ _17860_/Q _17861_/Q _12192_/C vssd1 vssd1 vccd1 vccd1 _12194_/B sky130_fd_sc_hd__and3_1
XFILLER_181_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11143_ _11143_/A1 _11141_/Y _11142_/X vssd1 vssd1 vccd1 vccd1 _11143_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_132_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19534_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15951_ _08825_/A _11977_/B _15955_/B _15854_/Y _16048_/A vssd1 vssd1 vccd1 vccd1
+ _15951_/X sky130_fd_sc_hd__a41o_1
X_11074_ _11568_/A _11072_/X _11073_/X _11570_/B1 vssd1 vssd1 vccd1 vccd1 _11074_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput120 dout1[21] vssd1 vssd1 vccd1 vccd1 input120/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput131 dout1[31] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_hd__clkbuf_2
XFILLER_209_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput142 dout1[41] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_hd__clkbuf_2
XFILLER_209_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10025_ _17895_/Q _15120_/A vssd1 vssd1 vccd1 vccd1 _10025_/Y sky130_fd_sc_hd__nor2_1
X_14902_ _15003_/A1 _13636_/Y _15003_/B1 _18647_/Q _15003_/C1 vssd1 vssd1 vccd1 vccd1
+ _14902_/X sky130_fd_sc_hd__a221o_1
Xinput153 dout1[51] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_hd__buf_2
X_18670_ _18715_/CLK _18670_/D vssd1 vssd1 vccd1 vccd1 _18670_/Q sky130_fd_sc_hd__dfxtp_1
X_15882_ _18669_/Q _15906_/A2 _15906_/B1 _15881_/X vssd1 vssd1 vccd1 vccd1 _15882_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput164 dout1[61] vssd1 vssd1 vccd1 vccd1 input164/X sky130_fd_sc_hd__buf_2
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 irq[13] vssd1 vssd1 vccd1 vccd1 input175/X sky130_fd_sc_hd__buf_2
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 irq[9] vssd1 vssd1 vccd1 vccd1 _15090_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17621_ _19488_/Q _15101_/A _17556_/A _17211_/B _17556_/X vssd1 vssd1 vccd1 vccd1
+ _17621_/X sky130_fd_sc_hd__a221o_1
Xinput197 localMemory_wb_adr_i[16] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__clkbuf_2
X_14833_ _15006_/A1 _14832_/X _14875_/B1 vssd1 vssd1 vccd1 vccd1 _14833_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ input104/X input75/X _14784_/S vssd1 vssd1 vccd1 vccd1 _14764_/X sky130_fd_sc_hd__mux2_8
X_17552_ _14268_/A _17528_/B _17214_/A _17551_/Y vssd1 vssd1 vccd1 vccd1 _17552_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _18737_/Q _18736_/Q _11976_/C vssd1 vssd1 vccd1 vccd1 _11977_/B sky130_fd_sc_hd__and3_1
XFILLER_263_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16503_ _17669_/A0 _19109_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _19109_/D sky130_fd_sc_hd__mux2_1
X_13715_ _17879_/Q _13747_/A2 _13714_/X _13747_/B2 vssd1 vssd1 vccd1 vccd1 _13715_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10927_ _10785_/A _10925_/X _10926_/X _11563_/B1 vssd1 vssd1 vccd1 vccd1 _10927_/X
+ sky130_fd_sc_hd__o31a_1
X_17483_ _17483_/A _17523_/B vssd1 vssd1 vccd1 vccd1 _17483_/Y sky130_fd_sc_hd__nand2_1
X_14695_ _16821_/A _14685_/X _14691_/X _14875_/A1 vssd1 vssd1 vccd1 vccd1 _14695_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19222_ _19623_/CLK _19222_/D vssd1 vssd1 vccd1 vccd1 _19222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16434_ _19042_/Q _17666_/A0 _16457_/S vssd1 vssd1 vccd1 vccd1 _19042_/D sky130_fd_sc_hd__mux2_1
X_13646_ _17941_/Q _13973_/A2 _13644_/Y _13645_/X _14342_/A vssd1 vssd1 vccd1 vccd1
+ _17941_/D sky130_fd_sc_hd__o221a_1
XFILLER_177_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10858_ _11584_/C1 _10855_/X _10857_/X vssd1 vssd1 vccd1 vccd1 _10858_/X sky130_fd_sc_hd__a21o_1
XFILLER_204_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16365_ _16465_/A0 _18976_/Q _16385_/S vssd1 vssd1 vccd1 vccd1 _18976_/D sky130_fd_sc_hd__mux2_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ _19602_/CLK _19153_/D vssd1 vssd1 vccd1 vccd1 _19153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _15452_/A _13574_/X _13576_/A _13970_/B2 vssd1 vssd1 vccd1 vccd1 _13577_/X
+ sky130_fd_sc_hd__a22o_1
X_10789_ _11579_/A _10767_/X _09107_/D vssd1 vssd1 vccd1 vccd1 _10789_/X sky130_fd_sc_hd__a21o_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18104_ _18734_/CLK _18104_/D vssd1 vssd1 vccd1 vccd1 _18104_/Q sky130_fd_sc_hd__dfxtp_4
X_15316_ _15342_/B _15315_/Y _15731_/B1 vssd1 vssd1 vccd1 vccd1 _15316_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12528_ _12577_/A _12538_/A _12528_/C _12514_/B vssd1 vssd1 vccd1 vccd1 _13165_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_8_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19084_ _19118_/CLK _19084_/D vssd1 vssd1 vccd1 vccd1 _19084_/Q sky130_fd_sc_hd__dfxtp_1
X_16296_ _17694_/A0 _18909_/Q _16325_/S vssd1 vssd1 vccd1 vccd1 _18909_/D sky130_fd_sc_hd__mux2_1
XFILLER_184_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18035_ _19573_/CLK _18035_/D vssd1 vssd1 vccd1 vccd1 _18035_/Q sky130_fd_sc_hd__dfxtp_1
X_15247_ _15271_/B _15247_/B vssd1 vssd1 vccd1 vccd1 _15250_/B sky130_fd_sc_hd__nor2_1
X_12459_ _14669_/B _16819_/C vssd1 vssd1 vccd1 vccd1 _12459_/X sky130_fd_sc_hd__or2_2
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15178_ _15179_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15200_/B sky130_fd_sc_hd__nor2_2
XFILLER_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14129_ _14510_/A0 _18068_/Q _14140_/S vssd1 vssd1 vccd1 vccd1 _18068_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18937_ _19648_/CLK _18937_/D vssd1 vssd1 vccd1 vccd1 _18937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_255_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09670_ _09690_/A _09665_/Y _09669_/Y _08843_/A vssd1 vssd1 vccd1 vccd1 _09670_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_95_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18868_ _19643_/CLK _18868_/D vssd1 vssd1 vccd1 vccd1 _18868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_283_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17819_ _19490_/CLK _17819_/D vssd1 vssd1 vccd1 vccd1 _17819_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18799_ _19607_/CLK _18799_/D vssd1 vssd1 vccd1 vccd1 _18799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09104_ _08948_/A _08948_/B _09102_/X vssd1 vssd1 vccd1 vccd1 _09104_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09035_ input117/X input153/X _09657_/S vssd1 vssd1 vccd1 vccd1 _09035_/X sky130_fd_sc_hd__mux2_8
XFILLER_163_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1808 _14442_/B vssd1 vssd1 vccd1 vccd1 _14449_/B sky130_fd_sc_hd__clkbuf_2
Xfanout810 _14454_/Y vssd1 vssd1 vccd1 vccd1 _14477_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_117_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout821 _14277_/S vssd1 vssd1 vccd1 vccd1 _14305_/S sky130_fd_sc_hd__clkbuf_16
Xfanout1819 _17380_/A vssd1 vssd1 vccd1 vccd1 _17366_/A sky130_fd_sc_hd__clkbuf_4
X_09937_ _18440_/Q _18341_/Q _09937_/S vssd1 vssd1 vccd1 vccd1 _09937_/X sky130_fd_sc_hd__mux2_1
Xfanout832 _16476_/A0 vssd1 vssd1 vccd1 vccd1 _16542_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout843 _17711_/A0 vssd1 vssd1 vccd1 vccd1 _17678_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_219_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout854 _10760_/X vssd1 vssd1 vccd1 vccd1 _10792_/A2 sky130_fd_sc_hd__buf_6
Xfanout865 _10341_/A2 vssd1 vssd1 vccd1 vccd1 _17719_/A0 sky130_fd_sc_hd__clkbuf_2
Xfanout876 _10166_/X vssd1 vssd1 vccd1 vccd1 _17721_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout887 _12935_/S vssd1 vssd1 vccd1 vccd1 _12943_/S sky130_fd_sc_hd__buf_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _08901_/A _19197_/Q _19165_/Q _09885_/S _08895_/A vssd1 vssd1 vccd1 vccd1
+ _09868_/X sky130_fd_sc_hd__a221o_1
Xfanout898 _17667_/A0 vssd1 vssd1 vccd1 vccd1 _16501_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _19448_/Q vssd1 vssd1 vccd1 vccd1 _08819_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09797_/X _09798_/X _11282_/A vssd1 vssd1 vccd1 vccd1 _09799_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_203 _14164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ _11865_/A _11828_/X _11829_/Y _11859_/B vssd1 vssd1 vccd1 vccd1 _11831_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _17906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_225 _18385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _18393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _18731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_258 input215/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _18579_/Q _14349_/B _11770_/B1 _13512_/B vssd1 vssd1 vccd1 vccd1 _11761_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 input230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _19441_/Q _13655_/A2 _13498_/X _13499_/X _13655_/C1 vssd1 vssd1 vccd1 vccd1
+ _13500_/X sky130_fd_sc_hd__o221a_1
XFILLER_242_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10703_/Y _10710_/Y _10711_/X _10697_/X vssd1 vssd1 vccd1 vccd1 _10712_/X
+ sky130_fd_sc_hd__o2bb2a_2
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _18332_/Q _16551_/A0 _14486_/S vssd1 vssd1 vccd1 vccd1 _18332_/D sky130_fd_sc_hd__mux2_1
X_11692_ _11692_/A1 _11690_/Y _11691_/X vssd1 vssd1 vccd1 vccd1 _11692_/X sky130_fd_sc_hd__o21a_2
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _19439_/Q _13655_/A2 _13429_/X _13430_/X _13655_/C1 vssd1 vssd1 vccd1 vccd1
+ _13431_/X sky130_fd_sc_hd__o221a_1
XFILLER_201_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10643_ _10641_/X _10642_/X _10643_/S vssd1 vssd1 vccd1 vccd1 _10643_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16150_ _16143_/C _18725_/Q _16141_/B vssd1 vssd1 vccd1 vccd1 _16150_/X sky130_fd_sc_hd__a21o_1
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13362_ _18114_/Q _13397_/C vssd1 vssd1 vccd1 vccd1 _13363_/A sky130_fd_sc_hd__xnor2_2
XFILLER_210_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10574_ _10649_/A1 _10573_/X _10572_/X _10881_/S1 vssd1 vssd1 vccd1 vccd1 _10574_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_182_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15101_ _15101_/A _15101_/B _15101_/C _15101_/D vssd1 vssd1 vccd1 vccd1 _17591_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_166_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12313_ _12315_/B _12314_/B vssd1 vssd1 vccd1 vccd1 _15329_/B sky130_fd_sc_hd__nor2_4
X_16081_ _18743_/Q _16093_/B vssd1 vssd1 vccd1 vccd1 _16081_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13293_ _14342_/A _13293_/B vssd1 vssd1 vccd1 vccd1 _17931_/D sky130_fd_sc_hd__and2_1
XFILLER_155_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15032_ _18521_/Q input198/X _15038_/S vssd1 vssd1 vccd1 vccd1 _18521_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12244_ _17880_/Q _12242_/B _12243_/Y vssd1 vssd1 vccd1 vccd1 _17880_/D sky130_fd_sc_hd__o21a_1
X_12175_ _17854_/Q _12176_/C _17855_/Q vssd1 vssd1 vccd1 vccd1 _12177_/B sky130_fd_sc_hd__a21oi_1
XFILLER_218_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11126_ _11352_/A1 _18324_/Q _17775_/Q _11353_/B2 vssd1 vssd1 vccd1 vccd1 _11126_/X
+ sky130_fd_sc_hd__a22o_1
X_16983_ _19328_/Q _17043_/B vssd1 vssd1 vccd1 vccd1 _16983_/X sky130_fd_sc_hd__or2_1
XFILLER_150_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18722_ _18772_/CLK _18722_/D vssd1 vssd1 vccd1 vccd1 _18722_/Q sky130_fd_sc_hd__dfxtp_1
X_15934_ _18687_/Q _15943_/A2 _15933_/X _15946_/C1 vssd1 vssd1 vccd1 vccd1 _18687_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_249_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ _18119_/Q _15502_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11061_/B sky130_fd_sc_hd__mux2_4
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10008_ _10707_/A _09997_/X _09998_/X _10007_/X _11237_/B1 vssd1 vssd1 vccd1 vccd1
+ _10009_/C sky130_fd_sc_hd__o311a_1
X_18653_ _19142_/CLK _18653_/D vssd1 vssd1 vccd1 vccd1 _18653_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15865_ _18664_/Q _15910_/A2 _15863_/X _15864_/X _15910_/C1 vssd1 vssd1 vccd1 vccd1
+ _18664_/D sky130_fd_sc_hd__o221a_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _19543_/Q _17622_/A2 _17591_/X _17184_/B _17603_/X vssd1 vssd1 vccd1 vccd1
+ _19543_/D sky130_fd_sc_hd__o221a_1
XFILLER_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14816_ _14696_/A _18270_/Q _14815_/Y _14918_/B1 vssd1 vssd1 vccd1 vccd1 _14816_/X
+ sky130_fd_sc_hd__a31o_2
X_18584_ _19481_/CLK _18584_/D vssd1 vssd1 vccd1 vccd1 _18584_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_184_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _19421_/Q _15796_/B vssd1 vssd1 vccd1 vccd1 _15796_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_92_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ _08883_/A _17532_/X _17533_/Y _17534_/X vssd1 vssd1 vccd1 vccd1 _17535_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14747_ _14718_/A _14746_/X _14846_/B1 vssd1 vssd1 vccd1 vccd1 _14747_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_33_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11959_ _19230_/Q _11959_/A2 _14345_/C _11959_/B2 vssd1 vssd1 vccd1 vccd1 _11959_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17466_ _18577_/Q _17527_/A1 _17516_/C1 vssd1 vssd1 vccd1 vccd1 _17466_/X sky130_fd_sc_hd__o21a_1
X_14678_ _14912_/A1 _12550_/X _14677_/X _18626_/Q _14973_/C1 vssd1 vssd1 vccd1 vccd1
+ _14678_/X sky130_fd_sc_hd__a221o_1
XFILLER_220_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19205_ _19594_/CLK _19205_/D vssd1 vssd1 vccd1 vccd1 _19205_/Q sky130_fd_sc_hd__dfxtp_1
X_16417_ _16615_/A0 _19026_/Q _16420_/S vssd1 vssd1 vccd1 vccd1 _19026_/D sky130_fd_sc_hd__mux2_1
X_13629_ _19511_/Q _13781_/A2 _13781_/B1 _13628_/X vssd1 vssd1 vccd1 vccd1 _13629_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17397_ _14423_/A _17396_/X _17437_/A2 _18778_/Q vssd1 vssd1 vccd1 vccd1 _17397_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19136_ _19608_/CLK _19136_/D vssd1 vssd1 vccd1 vccd1 _19136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16348_ _18960_/Q _17680_/A0 _16358_/S vssd1 vssd1 vccd1 vccd1 _18960_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16279_ _16610_/A0 _18893_/Q _16288_/S vssd1 vssd1 vccd1 vccd1 _18893_/D sky130_fd_sc_hd__mux2_1
X_19067_ _19195_/CLK _19067_/D vssd1 vssd1 vccd1 vccd1 _19067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput402 _11924_/X vssd1 vssd1 vccd1 vccd1 din0[4] sky130_fd_sc_hd__buf_4
X_18018_ _18973_/CLK _18018_/D vssd1 vssd1 vccd1 vccd1 _18018_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput413 _18483_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[12] sky130_fd_sc_hd__buf_4
Xoutput424 _18493_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[22] sky130_fd_sc_hd__buf_4
Xoutput435 _18474_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[3] sky130_fd_sc_hd__buf_4
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput446 _18734_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[1] sky130_fd_sc_hd__buf_4
Xoutput457 _14238_/A vssd1 vssd1 vccd1 vccd1 probe_programCounter[16] sky130_fd_sc_hd__buf_4
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput468 _18127_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[26] sky130_fd_sc_hd__buf_4
Xoutput479 _18108_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[7] sky130_fd_sc_hd__buf_4
XFILLER_271_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09722_ _19103_/Q _19135_/Q _09952_/S vssd1 vssd1 vccd1 vccd1 _09722_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09653_ _09992_/A _09653_/B vssd1 vssd1 vccd1 vccd1 _09653_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09584_ _09580_/X _09581_/X _10371_/S vssd1 vssd1 vccd1 vccd1 _09585_/B sky130_fd_sc_hd__mux2_1
XFILLER_270_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09018_ _09031_/S _09006_/X _09016_/X _08995_/B vssd1 vssd1 vccd1 vccd1 _09025_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_164_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10290_ _18622_/Q _18193_/Q _10290_/S vssd1 vssd1 vccd1 vccd1 _10290_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1605 _15104_/X vssd1 vssd1 vccd1 vccd1 _15116_/B sky130_fd_sc_hd__buf_4
XFILLER_132_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1616 _11141_/A vssd1 vssd1 vccd1 vccd1 _11556_/C sky130_fd_sc_hd__clkbuf_8
Xfanout1627 _09650_/B1 vssd1 vssd1 vccd1 vccd1 _09908_/B1 sky130_fd_sc_hd__buf_4
XFILLER_265_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1638 _09012_/A vssd1 vssd1 vccd1 vccd1 _11691_/B1 sky130_fd_sc_hd__buf_4
Xfanout640 _17345_/S vssd1 vssd1 vccd1 vccd1 _17377_/S sky130_fd_sc_hd__buf_6
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1649 _08901_/A vssd1 vssd1 vccd1 vccd1 _11618_/A1 sky130_fd_sc_hd__buf_8
Xfanout651 _17003_/B vssd1 vssd1 vccd1 vccd1 _17045_/B sky130_fd_sc_hd__buf_4
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout662 _13064_/B vssd1 vssd1 vccd1 vccd1 _13781_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_247_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13980_ _14004_/A _13980_/B vssd1 vssd1 vccd1 vccd1 _13980_/Y sky130_fd_sc_hd__nand2_1
XFILLER_282_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout673 _14996_/A1 vssd1 vssd1 vccd1 vccd1 _14875_/A1 sky130_fd_sc_hd__buf_4
XFILLER_247_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout684 _12564_/Y vssd1 vssd1 vccd1 vccd1 _12570_/C sky130_fd_sc_hd__buf_6
XFILLER_59_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout695 _13246_/A2 vssd1 vssd1 vccd1 vccd1 _13950_/A2 sky130_fd_sc_hd__buf_4
X_12931_ _12749_/X _12930_/X _13134_/S vssd1 vssd1 vccd1 vccd1 _12932_/B sky130_fd_sc_hd__mux2_2
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _17857_/Q _12919_/A2 _12850_/X _13303_/B2 _12861_/X vssd1 vssd1 vccd1 vccd1
+ _12862_/X sky130_fd_sc_hd__a221o_1
XFILLER_248_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15650_ _19480_/Q _19414_/Q vssd1 vssd1 vccd1 vccd1 _15651_/B sky130_fd_sc_hd__or2_1
XFILLER_74_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _16593_/A0 _18408_/Q _14630_/S vssd1 vssd1 vccd1 vccd1 _18408_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11813_ _11859_/A _11812_/X _11811_/Y vssd1 vssd1 vccd1 vccd1 _11814_/C sky130_fd_sc_hd__a21oi_4
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15581_ _18583_/Q _18582_/Q _15581_/C vssd1 vssd1 vccd1 vccd1 _15621_/C sky130_fd_sc_hd__and3_2
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _12672_/Y _12694_/X _12818_/S vssd1 vssd1 vccd1 vccd1 _12793_/X sky130_fd_sc_hd__mux2_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17320_ _17328_/A _17320_/B vssd1 vssd1 vccd1 vccd1 _19457_/D sky130_fd_sc_hd__and2_1
XFILLER_144_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14596_/A _14532_/B vssd1 vssd1 vccd1 vccd1 _18374_/D sky130_fd_sc_hd__or2_1
XFILLER_242_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11744_ _18568_/Q _14522_/A2 _11799_/B _13081_/A vssd1 vssd1 vccd1 vccd1 _11744_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _18315_/Q _16501_/A0 _14485_/S vssd1 vssd1 vccd1 vccd1 _18315_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17251_ _18111_/Q _17389_/B1 _17241_/B _19434_/Q vssd1 vssd1 vccd1 vccd1 _17251_/X
+ sky130_fd_sc_hd__a22o_1
X_11675_ _12593_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _13545_/B sky130_fd_sc_hd__xnor2_4
XFILLER_230_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16202_ _17699_/A0 _18818_/Q _16222_/S vssd1 vssd1 vccd1 vccd1 _18818_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ _13414_/A _13414_/B vssd1 vssd1 vccd1 vccd1 _13414_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17182_ _19412_/Q fanout533/X _17493_/A _17119_/B vssd1 vssd1 vccd1 vccd1 _17183_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_10626_ _11312_/A1 _17781_/Q _09108_/B _18330_/Q vssd1 vssd1 vccd1 vccd1 _10626_/X
+ sky130_fd_sc_hd__o22a_1
X_14394_ _16204_/A0 _18245_/Q _14415_/S vssd1 vssd1 vccd1 vccd1 _18245_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16133_ _18769_/Q _16141_/B vssd1 vssd1 vccd1 vccd1 _16133_/Y sky130_fd_sc_hd__nand2_1
XFILLER_167_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ _13928_/A1 _13334_/X _13344_/X vssd1 vssd1 vccd1 vccd1 _14000_/B sky130_fd_sc_hd__a21oi_4
XFILLER_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10557_ _10555_/X _10556_/X _10557_/S vssd1 vssd1 vccd1 vccd1 _10558_/B sky130_fd_sc_hd__mux2_1
XFILLER_170_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16064_ _16054_/A _16063_/B _16057_/X _16075_/A vssd1 vssd1 vccd1 vccd1 _16064_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13276_ _19243_/Q _13425_/A2 _13425_/B1 _19275_/Q vssd1 vssd1 vccd1 vccd1 _13276_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10488_ _10532_/A _17684_/A0 _10487_/Y _11800_/B vssd1 vssd1 vccd1 vccd1 _10489_/B
+ sky130_fd_sc_hd__o211ai_4
X_15015_ _18504_/Q input190/X _16627_/S vssd1 vssd1 vccd1 vccd1 _18504_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12227_ _12241_/A _12232_/C vssd1 vssd1 vccd1 vccd1 _12227_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12158_ _17848_/Q _12160_/C _12157_/Y vssd1 vssd1 vccd1 vccd1 _17848_/D sky130_fd_sc_hd__o21a_1
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11109_ _11107_/X _11108_/X _11127_/S vssd1 vssd1 vccd1 vccd1 _11109_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16966_ _16970_/A1 _17950_/Q _16965_/X vssd1 vssd1 vccd1 vccd1 _17211_/B sky130_fd_sc_hd__o21a_4
X_12089_ _12089_/A _14224_/B vssd1 vssd1 vccd1 vccd1 _12089_/Y sky130_fd_sc_hd__nand2_1
XFILLER_238_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18705_ _19306_/CLK _18705_/D vssd1 vssd1 vccd1 vccd1 _18705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15917_ _15917_/A _15941_/S _15923_/C vssd1 vssd1 vccd1 vccd1 _15917_/X sky130_fd_sc_hd__and3_1
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16897_ _18755_/Q _16961_/A2 _16969_/B1 input219/X _08828_/A vssd1 vssd1 vccd1 vccd1
+ _16897_/X sky130_fd_sc_hd__a221o_1
XFILLER_265_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18636_ _19142_/CLK _18636_/D vssd1 vssd1 vccd1 vccd1 _18636_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_225_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _16041_/A _16063_/A vssd1 vssd1 vccd1 vccd1 _15854_/B sky130_fd_sc_hd__or2_4
XFILLER_264_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18567_ _19525_/CLK _18567_/D vssd1 vssd1 vccd1 vccd1 _18567_/Q sky130_fd_sc_hd__dfxtp_4
X_15779_ _15753_/Y _15758_/B _15755_/B vssd1 vssd1 vccd1 vccd1 _15780_/B sky130_fd_sc_hd__o21ai_2
XFILLER_80_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17518_ _18126_/Q _17528_/B _17516_/X _17517_/Y vssd1 vssd1 vccd1 vccd1 _17518_/X
+ sky130_fd_sc_hd__a211o_1
X_18498_ _18501_/CLK _18498_/D vssd1 vssd1 vccd1 vccd1 _18498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17449_ _19501_/Q _17453_/B _17447_/X _17448_/Y _17326_/A vssd1 vssd1 vccd1 vccd1
+ _19501_/D sky130_fd_sc_hd__o221a_1
XFILLER_220_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19119_ _19618_/CLK _19119_/D vssd1 vssd1 vccd1 vccd1 _19119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput287 _11962_/X vssd1 vssd1 vccd1 vccd1 addr0[2] sky130_fd_sc_hd__buf_4
Xoutput298 _11914_/X vssd1 vssd1 vccd1 vccd1 addr1[4] sky130_fd_sc_hd__buf_4
XFILLER_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09705_ _10366_/A1 _19199_/Q _19167_/Q _09720_/S _12766_/A0 vssd1 vssd1 vccd1 vccd1
+ _09705_/X sky130_fd_sc_hd__a221o_1
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09636_ _18444_/Q _18345_/Q _10313_/S vssd1 vssd1 vccd1 vccd1 _09636_/X sky130_fd_sc_hd__mux2_1
XFILLER_215_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09567_ _09992_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09567_/Y sky130_fd_sc_hd__nand2_1
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09498_ _18600_/Q _18171_/Q _09498_/S vssd1 vssd1 vccd1 vccd1 _09498_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ _18544_/Q _11462_/S vssd1 vssd1 vccd1 vccd1 _11460_/X sky130_fd_sc_hd__or2_1
XFILLER_109_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10411_ _09135_/S _10410_/X _11459_/B1 vssd1 vssd1 vccd1 vccd1 _10411_/X sky130_fd_sc_hd__o21a_1
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ _18452_/Q _18353_/Q _11477_/S vssd1 vssd1 vccd1 vccd1 _11391_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13130_ _13130_/A _13130_/B vssd1 vssd1 vccd1 vccd1 _13130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10342_ _11411_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10342_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13061_ _19238_/Q _13495_/A2 _13495_/B1 _19270_/Q vssd1 vssd1 vccd1 vccd1 _13061_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10273_ _18335_/Q _17786_/Q _10299_/S vssd1 vssd1 vccd1 vccd1 _10273_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12012_ _17779_/Q _17680_/A0 _12022_/S vssd1 vssd1 vccd1 vccd1 _17779_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1402 _09542_/S vssd1 vssd1 vccd1 vccd1 _09680_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1413 fanout1415/X vssd1 vssd1 vccd1 vccd1 _09181_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_279_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1424 _11403_/S vssd1 vssd1 vccd1 vccd1 _11455_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_39_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19622_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16820_ _16821_/A _12461_/A _16820_/A3 _16819_/Y vssd1 vssd1 vccd1 vccd1 _16839_/B
+ sky130_fd_sc_hd__a31o_1
Xfanout1435 _10557_/S vssd1 vssd1 vccd1 vccd1 _11562_/S sky130_fd_sc_hd__buf_6
Xfanout1446 _09087_/Y vssd1 vssd1 vccd1 vccd1 _11002_/C1 sky130_fd_sc_hd__buf_6
Xfanout1457 _09086_/Y vssd1 vssd1 vccd1 vccd1 _10337_/S1 sky130_fd_sc_hd__buf_12
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1468 fanout1469/X vssd1 vssd1 vccd1 vccd1 _11605_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_266_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1479 _09801_/S vssd1 vssd1 vccd1 vccd1 _11609_/S sky130_fd_sc_hd__buf_4
X_16751_ _19270_/Q _19269_/Q _16751_/C vssd1 vssd1 vccd1 vccd1 _16754_/B sky130_fd_sc_hd__and3_1
Xfanout492 _14667_/X vssd1 vssd1 vccd1 vccd1 _14889_/B1 sky130_fd_sc_hd__clkbuf_16
XFILLER_247_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13963_ _13962_/A _12756_/Y _13962_/B vssd1 vssd1 vccd1 vccd1 _13963_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15702_ _15702_/A _15702_/B vssd1 vssd1 vccd1 vccd1 _15707_/A sky130_fd_sc_hd__xnor2_2
XFILLER_111_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12914_ _19363_/Q _12913_/X _13925_/S vssd1 vssd1 vccd1 vccd1 _12914_/X sky130_fd_sc_hd__mux2_2
X_19470_ _19470_/CLK _19470_/D vssd1 vssd1 vccd1 vccd1 _19470_/Q sky130_fd_sc_hd__dfxtp_2
X_16682_ _19247_/Q _19243_/Q _19239_/Q _19234_/Q vssd1 vssd1 vccd1 vccd1 _16683_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_207_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13894_ _11634_/B _13912_/A2 _14153_/A vssd1 vssd1 vccd1 vccd1 _13894_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_262_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18421_ _18613_/CLK _18421_/D vssd1 vssd1 vccd1 vccd1 _18421_/Q sky130_fd_sc_hd__dfxtp_1
X_15633_ _15625_/Y _15626_/X _15632_/X _15717_/B2 _15633_/C1 vssd1 vssd1 vccd1 vccd1
+ _15633_/X sky130_fd_sc_hd__a221o_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ _09948_/X _13292_/A2 _12844_/X _13256_/B1 _17921_/Q vssd1 vssd1 vccd1 vccd1
+ _12846_/B sky130_fd_sc_hd__a32o_1
XFILLER_234_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _19208_/CLK _18352_/D vssd1 vssd1 vccd1 vccd1 _18352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _19361_/Q _12775_/X _13925_/S vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__mux2_2
X_15564_ _19444_/Q _15793_/A2 _17208_/A vssd1 vssd1 vccd1 vccd1 _15564_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17303_ _17301_/Y _17302_/X _17198_/A vssd1 vssd1 vccd1 vccd1 _19451_/D sky130_fd_sc_hd__a21oi_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14515_ _17717_/A0 _18365_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _18365_/D sky130_fd_sc_hd__mux2_1
X_11727_ _17531_/A _11727_/B vssd1 vssd1 vccd1 vccd1 _11728_/C sky130_fd_sc_hd__nor2_1
X_18283_ _19448_/CLK _18283_/D vssd1 vssd1 vccd1 vccd1 _18283_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _19473_/Q _19407_/Q vssd1 vssd1 vccd1 vccd1 _15496_/B sky130_fd_sc_hd__or2_2
XFILLER_203_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17234_ _17232_/Y _17233_/X _14423_/B vssd1 vssd1 vccd1 vccd1 _19428_/D sky130_fd_sc_hd__a21oi_1
X_14446_ _18585_/Q _17376_/A vssd1 vssd1 vccd1 vccd1 _18298_/D sky130_fd_sc_hd__and2_1
X_11658_ _15082_/B _12837_/B vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__nand2_8
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10609_ _17943_/Q _08948_/B _10608_/X vssd1 vssd1 vccd1 vccd1 _10609_/X sky130_fd_sc_hd__o21a_4
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14377_ _18229_/Q _16551_/A0 _14377_/S vssd1 vssd1 vccd1 vccd1 _18229_/D sky130_fd_sc_hd__mux2_1
X_17165_ _17231_/A _17165_/B vssd1 vssd1 vccd1 vccd1 _19406_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11589_ _09107_/D _11579_/Y _11588_/Y _09859_/A vssd1 vssd1 vccd1 vccd1 _11589_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_128_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16116_ _16140_/A1 _16115_/Y _16142_/B1 vssd1 vssd1 vccd1 vccd1 _18760_/D sky130_fd_sc_hd__a21oi_1
XFILLER_143_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13328_ _15382_/B2 _13324_/X _13327_/X _13936_/B2 vssd1 vssd1 vccd1 vccd1 _13329_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17096_ _17184_/B _17108_/A2 _17095_/X _17360_/A vssd1 vssd1 vccd1 vccd1 _19381_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16047_ _18728_/Q _18735_/Q _16051_/S vssd1 vssd1 vccd1 vccd1 _16048_/B sky130_fd_sc_hd__mux2_1
X_13259_ _13260_/A _13260_/B vssd1 vssd1 vccd1 vccd1 _13259_/X sky130_fd_sc_hd__and2_4
XFILLER_89_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17998_ _18613_/CLK _17998_/D vssd1 vssd1 vccd1 vccd1 _17998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16949_ _18768_/Q _16965_/A2 _16965_/B1 input233/X _16965_/C1 vssd1 vssd1 vccd1 vccd1
+ _16949_/X sky130_fd_sc_hd__a221o_2
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09421_ _10294_/A1 _19106_/Q _19138_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09421_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18619_ _19643_/CLK _18619_/D vssd1 vssd1 vccd1 vccd1 _18619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19599_ _19599_/CLK _19599_/D vssd1 vssd1 vccd1 vccd1 _19599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _09350_/X _09351_/X _10409_/A vssd1 vssd1 vccd1 vccd1 _09352_/X sky130_fd_sc_hd__mux2_1
XFILLER_212_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09283_ _11498_/A1 _18142_/Q _18788_/Q _09302_/S _10144_/B1 vssd1 vssd1 vccd1 vccd1
+ _09283_/X sky130_fd_sc_hd__a221o_1
XFILLER_221_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ _09245_/A _11556_/A _11556_/B _08997_/X vssd1 vssd1 vccd1 vccd1 _11218_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10960_ _11352_/A1 _19118_/Q _19150_/Q _11125_/B2 vssd1 vssd1 vccd1 vccd1 _10960_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _10323_/A1 _19136_/Q _11171_/S _19104_/Q vssd1 vssd1 vccd1 vccd1 _09619_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10891_ _18863_/Q _18895_/Q _19055_/Q _19023_/Q _10815_/B _11357_/S1 vssd1 vssd1
+ vccd1 vccd1 _10891_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12630_ _13411_/A _12596_/Y _12629_/X _12595_/Y vssd1 vssd1 vccd1 vccd1 _13465_/C
+ sky130_fd_sc_hd__a211oi_4
Xclkbuf_leaf_157_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19477_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12561_ _12577_/A _12561_/B vssd1 vssd1 vccd1 vccd1 _12562_/B sky130_fd_sc_hd__or2_1
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11512_ _11512_/A1 _19630_/Q _18919_/Q _11513_/B2 vssd1 vssd1 vccd1 vccd1 _11512_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14300_ _17718_/A0 _18159_/Q _14305_/S vssd1 vssd1 vccd1 vccd1 _18159_/D sky130_fd_sc_hd__mux2_1
X_15280_ _15280_/A _15280_/B vssd1 vssd1 vccd1 vccd1 _15280_/X sky130_fd_sc_hd__xor2_1
X_12492_ _12492_/A _12492_/B vssd1 vssd1 vccd1 vccd1 _12492_/X sky130_fd_sc_hd__and2_2
XFILLER_157_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ _18287_/Q _14247_/A2 _14230_/X _15718_/C1 vssd1 vssd1 vccd1 vccd1 _18113_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11443_ _12597_/B vssd1 vssd1 vccd1 vccd1 _11445_/B sky130_fd_sc_hd__clkinv_2
XFILLER_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14162_ _18731_/Q _15954_/B vssd1 vssd1 vccd1 vccd1 _15953_/A sky130_fd_sc_hd__nand2_2
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11374_ _09987_/A _11373_/X _11371_/X vssd1 vssd1 vccd1 vccd1 _11374_/X sky130_fd_sc_hd__o21a_1
XFILLER_153_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13113_ input8/X _12552_/X _13106_/X _13112_/X _12538_/B vssd1 vssd1 vccd1 vccd1
+ _13113_/X sky130_fd_sc_hd__o221a_2
XFILLER_180_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10325_ _10315_/X _10318_/X _10321_/X _10324_/X _10689_/S _09350_/S vssd1 vssd1 vccd1
+ vccd1 _10326_/B sky130_fd_sc_hd__mux4_2
X_14093_ _16609_/A0 _18033_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _18033_/D sky130_fd_sc_hd__mux2_1
X_18970_ _19163_/CLK _18970_/D vssd1 vssd1 vccd1 vccd1 _18970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13044_ _13797_/A0 _12756_/Y _13044_/S vssd1 vssd1 vccd1 vccd1 _13044_/X sky130_fd_sc_hd__mux2_1
X_17921_ _17930_/CLK _17921_/D vssd1 vssd1 vccd1 vccd1 _17921_/Q sky130_fd_sc_hd__dfxtp_4
X_10256_ _18560_/Q _18435_/Q _18044_/Q _18012_/Q _10253_/C _10266_/S1 vssd1 vssd1
+ vccd1 vccd1 _10256_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1210 _14154_/B1 vssd1 vssd1 vccd1 vccd1 _12704_/S sky130_fd_sc_hd__buf_4
Xfanout1221 _13899_/A vssd1 vssd1 vccd1 vccd1 _15133_/A sky130_fd_sc_hd__buf_8
X_17852_ _19261_/CLK _17852_/D vssd1 vssd1 vccd1 vccd1 _17852_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1232 _12277_/Y vssd1 vssd1 vccd1 vccd1 _14692_/A2 sky130_fd_sc_hd__buf_4
XFILLER_120_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10187_ _10334_/A1 _18233_/Q _10090_/S _18968_/Q vssd1 vssd1 vccd1 vccd1 _10187_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1243 _09033_/X vssd1 vssd1 vccd1 vccd1 _09034_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_67_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1254 _10905_/S vssd1 vssd1 vccd1 vccd1 _13904_/A sky130_fd_sc_hd__buf_6
XFILLER_267_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16803_ _16803_/A _16803_/B _16807_/C vssd1 vssd1 vccd1 vccd1 _19289_/D sky130_fd_sc_hd__nor3_1
XFILLER_38_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1265 _09866_/B vssd1 vssd1 vccd1 vccd1 _09946_/B1 sky130_fd_sc_hd__buf_8
Xfanout1276 _14875_/B1 vssd1 vssd1 vccd1 vccd1 _14865_/B1 sky130_fd_sc_hd__buf_8
XFILLER_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1287 _15037_/S vssd1 vssd1 vccd1 vccd1 _16627_/S sky130_fd_sc_hd__buf_6
X_17783_ _19611_/CLK _17783_/D vssd1 vssd1 vccd1 vccd1 _17783_/Q sky130_fd_sc_hd__dfxtp_1
X_14995_ _14995_/A1 _14993_/X _14994_/X _14934_/X vssd1 vssd1 vccd1 vccd1 _14995_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1298 _14524_/X vssd1 vssd1 vccd1 vccd1 _14586_/A sky130_fd_sc_hd__buf_4
XFILLER_75_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19522_ _19522_/CLK _19522_/D vssd1 vssd1 vccd1 vccd1 _19522_/Q sky130_fd_sc_hd__dfxtp_1
X_16734_ _19264_/Q _19263_/Q _16734_/C vssd1 vssd1 vccd1 vccd1 _16739_/C sky130_fd_sc_hd__and3_1
X_13946_ _19553_/Q _13946_/B vssd1 vssd1 vccd1 vccd1 _13946_/X sky130_fd_sc_hd__or2_1
XFILLER_62_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19453_ _19453_/CLK _19453_/D vssd1 vssd1 vccd1 vccd1 _19453_/Q sky130_fd_sc_hd__dfxtp_1
X_16665_ _16768_/A _16665_/B _16670_/C vssd1 vssd1 vccd1 vccd1 _19243_/D sky130_fd_sc_hd__nor3_1
XFILLER_262_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13877_ _19261_/Q _13943_/A2 _13943_/B1 _19293_/Q vssd1 vssd1 vccd1 vccd1 _13877_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18404_ _19464_/CLK _18404_/D vssd1 vssd1 vccd1 vccd1 _18404_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15616_ _13679_/A _15111_/A _13706_/X _15112_/B vssd1 vssd1 vccd1 vccd1 _15616_/X
+ sky130_fd_sc_hd__o22a_1
X_12828_ _12817_/Y _12827_/X _13135_/S vssd1 vssd1 vccd1 vccd1 _12828_/X sky130_fd_sc_hd__mux2_2
XFILLER_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19384_ _19483_/CLK _19384_/D vssd1 vssd1 vccd1 vccd1 _19384_/Q sky130_fd_sc_hd__dfxtp_2
X_16596_ _17696_/A0 _19199_/Q _16619_/S vssd1 vssd1 vccd1 vccd1 _19199_/D sky130_fd_sc_hd__mux2_1
X_18335_ _19159_/CLK _18335_/D vssd1 vssd1 vccd1 vccd1 _18335_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _18581_/Q _15718_/A2 _15546_/X _17356_/A vssd1 vssd1 vccd1 vccd1 _18581_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _11859_/A _12837_/B _14155_/A _11647_/A vssd1 vssd1 vccd1 vccd1 _12759_/X
+ sky130_fd_sc_hd__o22a_1
X_18266_ _19628_/CLK _18266_/D vssd1 vssd1 vccd1 vccd1 _18266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15478_ _15478_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _15478_/Y sky130_fd_sc_hd__nor2_1
X_17217_ _17217_/A _17217_/B vssd1 vssd1 vccd1 vccd1 _17250_/B sky130_fd_sc_hd__or2_4
X_14429_ _18568_/Q _16052_/A vssd1 vssd1 vccd1 vccd1 _18281_/D sky130_fd_sc_hd__and2_1
X_18197_ _18817_/CLK _18197_/D vssd1 vssd1 vccd1 vccd1 _18197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17148_ _17166_/A _17577_/A vssd1 vssd1 vccd1 vccd1 _17438_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09970_ _18627_/Q _18049_/Q _09973_/S vssd1 vssd1 vccd1 vccd1 _09970_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17079_ _19373_/Q _17113_/B vssd1 vssd1 vccd1 vccd1 _17079_/X sky130_fd_sc_hd__or2_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08921_ _12089_/A _17797_/Q vssd1 vssd1 vccd1 vccd1 _16459_/A sky130_fd_sc_hd__and2_4
XFILLER_130_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08852_ _17898_/Q vssd1 vssd1 vccd1 vccd1 _08852_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ _13148_/A vssd1 vssd1 vccd1 vccd1 _09404_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09335_ _18141_/Q _18787_/Q _09937_/S vssd1 vssd1 vccd1 vccd1 _09335_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09266_ _09264_/X _09265_/X _10409_/A vssd1 vssd1 vccd1 vccd1 _09266_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09197_ _18246_/Q _18821_/Q _10128_/B vssd1 vssd1 vccd1 vccd1 _09197_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10110_ _10336_/A _10109_/X _11466_/B1 vssd1 vssd1 vccd1 vccd1 _10110_/X sky130_fd_sc_hd__o21a_1
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11090_ _18828_/Q _11300_/B vssd1 vssd1 vccd1 vccd1 _11090_/X sky130_fd_sc_hd__or2_1
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ _10589_/S _10041_/B vssd1 vssd1 vccd1 vccd1 _10041_/Y sky130_fd_sc_hd__nor2_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ _13966_/C1 _13799_/X _13796_/Y vssd1 vssd1 vccd1 vccd1 _13800_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11992_ _17759_/Q _16593_/A0 _12019_/S vssd1 vssd1 vccd1 vccd1 _17759_/D sky130_fd_sc_hd__mux2_1
X_14780_ _14992_/A1 _13217_/X _14973_/B1 _18635_/Q _14741_/B vssd1 vssd1 vccd1 vccd1
+ _14780_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13731_ _10604_/Y _13797_/A0 _13730_/Y _10603_/B vssd1 vssd1 vccd1 vccd1 _13731_/X
+ sky130_fd_sc_hd__o22a_1
X_10943_ _10937_/X _10939_/X _10942_/X _11578_/S _11588_/B1 vssd1 vssd1 vccd1 vccd1
+ _10943_/X sky130_fd_sc_hd__o221a_1
XFILLER_244_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16450_ _19058_/Q _16615_/A0 _16453_/S vssd1 vssd1 vccd1 vccd1 _19058_/D sky130_fd_sc_hd__mux2_1
X_13662_ _13931_/A _13660_/Y _13661_/X _13676_/B _13294_/A vssd1 vssd1 vccd1 vccd1
+ _13662_/X sky130_fd_sc_hd__o32a_1
X_10874_ _10027_/A _11135_/S _11181_/B1 _10873_/Y vssd1 vssd1 vccd1 vccd1 _12641_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15401_ _17129_/A _15400_/X _15499_/B1 vssd1 vssd1 vccd1 vccd1 _15401_/X sky130_fd_sc_hd__a21o_1
X_12613_ _09561_/B _12613_/B vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__nand2b_1
X_13593_ _13682_/B2 _13582_/X _13583_/Y _13592_/Y vssd1 vssd1 vccd1 vccd1 _14014_/B
+ sky130_fd_sc_hd__o2bb2a_4
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16381_ _16547_/A0 _18992_/Q _16391_/S vssd1 vssd1 vccd1 vccd1 _18992_/D sky130_fd_sc_hd__mux2_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18120_ _18741_/CLK _18120_/D vssd1 vssd1 vccd1 vccd1 _18120_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12544_ _12544_/A _12579_/A vssd1 vssd1 vccd1 vccd1 _12544_/Y sky130_fd_sc_hd__nor2_4
X_15332_ _15332_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15332_/X sky130_fd_sc_hd__and2_1
XFILLER_200_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18051_ _19114_/CLK _18051_/D vssd1 vssd1 vccd1 vccd1 _18051_/Q sky130_fd_sc_hd__dfxtp_1
X_12475_ _12488_/A _17916_/Q _12474_/Y vssd1 vssd1 vccd1 vccd1 _12501_/A sky130_fd_sc_hd__a21o_1
X_15263_ _15179_/B _15207_/A _15263_/C _15263_/D vssd1 vssd1 vccd1 vccd1 _15263_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17002_ _17577_/A _17032_/A2 _17001_/X _17469_/C1 vssd1 vssd1 vccd1 vccd1 _19337_/D
+ sky130_fd_sc_hd__o211a_1
X_11426_ _11506_/A1 _19112_/Q _19144_/Q _11426_/B2 vssd1 vssd1 vccd1 vccd1 _11426_/X
+ sky130_fd_sc_hd__a22o_1
X_14214_ _14214_/A _14244_/B vssd1 vssd1 vccd1 vccd1 _14214_/X sky130_fd_sc_hd__or2_1
XANTENNA_6 _18202_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ _15194_/A _15259_/B vssd1 vssd1 vccd1 vccd1 _15194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_54_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19193_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_153_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ _14145_/A _14145_/B _14145_/C vssd1 vssd1 vccd1 vccd1 _14146_/C sky130_fd_sc_hd__or3_1
X_11357_ _18250_/Q _18825_/Q _18453_/Q _18354_/Q _11360_/B2 _11357_/S1 vssd1 vssd1
+ vccd1 vccd1 _11358_/B sky130_fd_sc_hd__mux4_2
XFILLER_126_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10308_ _10308_/A vssd1 vssd1 vccd1 vccd1 _11636_/B sky130_fd_sc_hd__clkinv_2
XFILLER_152_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18953_ _19600_/CLK _18953_/D vssd1 vssd1 vccd1 vccd1 _18953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14076_ _17659_/A0 _18016_/Q _14098_/S vssd1 vssd1 vccd1 vccd1 _18016_/D sky130_fd_sc_hd__mux2_1
X_11288_ _11131_/A _11267_/Y _11273_/Y _11280_/Y _11287_/X vssd1 vssd1 vccd1 vccd1
+ _11288_/X sky130_fd_sc_hd__o32a_4
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17904_ _19595_/CLK _17904_/D vssd1 vssd1 vccd1 vccd1 _17904_/Q sky130_fd_sc_hd__dfxtp_4
X_13027_ _13462_/A _13027_/B _13027_/C vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__and3_1
X_10239_ _10239_/A _10239_/B vssd1 vssd1 vccd1 vccd1 _10239_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18884_ _18884_/CLK _18884_/D vssd1 vssd1 vccd1 vccd1 _18884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1040 _11411_/A vssd1 vssd1 vccd1 vccd1 _11488_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_266_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1051 _08883_/Y vssd1 vssd1 vccd1 vccd1 _17528_/B sky130_fd_sc_hd__buf_6
XFILLER_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17835_ _19300_/CLK _17835_/D vssd1 vssd1 vccd1 vccd1 _17835_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1062 _13958_/B vssd1 vssd1 vccd1 vccd1 _13761_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_66_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1073 _14027_/A2 vssd1 vssd1 vccd1 vccd1 _14032_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1084 _09911_/X vssd1 vssd1 vccd1 vccd1 _09980_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_281_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1095 _11210_/A1 vssd1 vssd1 vccd1 vccd1 _11518_/B2 sky130_fd_sc_hd__clkbuf_16
XFILLER_282_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17766_ _19126_/CLK _17766_/D vssd1 vssd1 vccd1 vccd1 _17766_/Q sky130_fd_sc_hd__dfxtp_1
X_14978_ _14978_/A vssd1 vssd1 vccd1 vccd1 _14978_/Y sky130_fd_sc_hd__clkinv_4
X_19505_ _19537_/CLK _19505_/D vssd1 vssd1 vccd1 vccd1 _19505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16717_ _19258_/Q _19257_/Q _19256_/Q _16717_/D vssd1 vssd1 vccd1 vccd1 _16723_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_63_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13929_ _13929_/A1 _13928_/X _13917_/Y vssd1 vssd1 vccd1 vccd1 _13931_/B sky130_fd_sc_hd__a21oi_1
X_17697_ _17697_/A0 _19623_/Q _17719_/S vssd1 vssd1 vccd1 vccd1 _19623_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19436_ _19464_/CLK _19436_/D vssd1 vssd1 vccd1 vccd1 _19436_/Q sky130_fd_sc_hd__dfxtp_2
X_16648_ _16648_/A _16648_/B vssd1 vssd1 vccd1 vccd1 _19238_/D sky130_fd_sc_hd__nor2_1
XFILLER_228_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19367_ _19464_/CLK _19367_/D vssd1 vssd1 vccd1 vccd1 _19367_/Q sky130_fd_sc_hd__dfxtp_1
X_16579_ _17712_/A0 _19183_/Q _16585_/S vssd1 vssd1 vccd1 vccd1 _19183_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09120_ _09117_/X _09119_/X _12408_/A vssd1 vssd1 vccd1 vccd1 _09120_/X sky130_fd_sc_hd__a21bo_1
X_18318_ _19565_/CLK _18318_/D vssd1 vssd1 vccd1 vccd1 _18318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19298_ _19326_/CLK _19298_/D vssd1 vssd1 vccd1 vccd1 _19298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09051_ _09030_/X _09038_/X _09047_/X _09050_/X vssd1 vssd1 vccd1 vccd1 _09052_/B
+ sky130_fd_sc_hd__o22a_1
X_18249_ _19075_/CLK _18249_/D vssd1 vssd1 vccd1 vccd1 _18249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09953_ _09951_/X _09952_/X _09972_/S vssd1 vssd1 vccd1 vccd1 _09953_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08904_ _08904_/A _09429_/S _08904_/C vssd1 vssd1 vccd1 vccd1 _08958_/A sky130_fd_sc_hd__and3_2
X_09884_ _18050_/Q _10816_/A2 _09883_/X _11189_/A vssd1 vssd1 vccd1 vccd1 _09884_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08835_ _18103_/Q vssd1 vssd1 vccd1 vccd1 _14714_/A sky130_fd_sc_hd__inv_6
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_407 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_418 _15357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_429 _11836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09318_ _13195_/S _09318_/B vssd1 vssd1 vccd1 vccd1 _13188_/A sky130_fd_sc_hd__nand2_2
X_10590_ _10663_/S _10583_/X _10584_/X vssd1 vssd1 vccd1 vccd1 _10590_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_278_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ _18142_/Q _18788_/Q _09252_/S vssd1 vssd1 vccd1 vccd1 _09249_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _17886_/Q _12257_/B _12259_/Y vssd1 vssd1 vccd1 vccd1 _17886_/D sky130_fd_sc_hd__o21a_1
XFILLER_181_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11211_ _14238_/A _15450_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11214_/B sky130_fd_sc_hd__mux2_4
XFILLER_123_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12191_ _17860_/Q _12192_/C _17861_/Q vssd1 vssd1 vccd1 vccd1 _12193_/B sky130_fd_sc_hd__a21oi_1
XFILLER_147_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11142_ _17968_/Q _11295_/A2 _11216_/B1 vssd1 vssd1 vccd1 vccd1 _11142_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15950_ _08825_/A _11977_/B _15849_/A _18693_/Q vssd1 vssd1 vccd1 vccd1 _15952_/B
+ sky130_fd_sc_hd__a31o_1
X_11073_ _11565_/A1 _19148_/Q _11073_/B1 _19116_/Q _11562_/S vssd1 vssd1 vccd1 vccd1
+ _11073_/X sky130_fd_sc_hd__o221a_1
XFILLER_277_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput110 dout1[12] vssd1 vssd1 vccd1 vccd1 input110/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput121 dout1[22] vssd1 vssd1 vccd1 vccd1 input121/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput132 dout1[32] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10024_ _11333_/A1 _17659_/A0 _10023_/X _11257_/C1 vssd1 vssd1 vccd1 vccd1 _11782_/B
+ sky130_fd_sc_hd__o211ai_4
X_14901_ _17811_/Q _15002_/B vssd1 vssd1 vccd1 vccd1 _14901_/X sky130_fd_sc_hd__or2_1
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput143 dout1[42] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput154 dout1[52] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_hd__buf_2
X_15881_ _15881_/A _15881_/B _15908_/C vssd1 vssd1 vccd1 vccd1 _15881_/X sky130_fd_sc_hd__and3_1
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput165 dout1[62] vssd1 vssd1 vccd1 vccd1 input165/X sky130_fd_sc_hd__buf_2
XFILLER_263_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 irq[14] vssd1 vssd1 vccd1 vccd1 _15087_/C sky130_fd_sc_hd__buf_4
X_17620_ _19551_/Q _17624_/A2 _17591_/X _17208_/B _17619_/X vssd1 vssd1 vccd1 vccd1
+ _19551_/D sky130_fd_sc_hd__o221a_1
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _14964_/B1 _14830_/X _14831_/X _14771_/X vssd1 vssd1 vccd1 vccd1 _14832_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_172_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19485_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput187 jtag_tck vssd1 vssd1 vccd1 vccd1 _16038_/A sky130_fd_sc_hd__buf_4
Xinput198 localMemory_wb_adr_i[17] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__clkbuf_2
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_101_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18666_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17551_ _18593_/Q _17538_/A _17550_/Y _17528_/B vssd1 vssd1 vccd1 vccd1 _17551_/Y
+ sky130_fd_sc_hd__a211oi_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14763_ _14865_/A1 _14762_/X _14865_/B1 vssd1 vssd1 vccd1 vccd1 _14763_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_251_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11975_ _18735_/Q _18734_/Q _18733_/Q vssd1 vssd1 vccd1 vccd1 _11976_/C sky130_fd_sc_hd__and3_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _16535_/A0 _19108_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _19108_/D sky130_fd_sc_hd__mux2_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13714_ _19256_/Q _13943_/A2 _13943_/B1 _19288_/Q vssd1 vssd1 vccd1 vccd1 _13714_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10926_ _11572_/A1 _17777_/Q _10940_/S _18326_/Q _10784_/S vssd1 vssd1 vccd1 vccd1
+ _10926_/X sky130_fd_sc_hd__o221a_1
X_17482_ _18119_/Q _17539_/C1 _17480_/X _17481_/X vssd1 vssd1 vccd1 vccd1 _17482_/X
+ sky130_fd_sc_hd__a22o_1
X_14694_ _16819_/B _14693_/Y _12277_/A vssd1 vssd1 vccd1 vccd1 _14694_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19221_ _19644_/CLK _19221_/D vssd1 vssd1 vccd1 vccd1 _19221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16433_ _19041_/Q _17665_/A0 _16454_/S vssd1 vssd1 vccd1 vccd1 _19041_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10857_ _19215_/Q _11482_/A2 _10856_/X _11578_/S vssd1 vssd1 vccd1 vccd1 _10857_/X
+ sky130_fd_sc_hd__a211o_1
X_13645_ _13938_/A _13622_/B _13971_/A2 _10471_/S _13579_/A vssd1 vssd1 vccd1 vccd1
+ _13645_/X sky130_fd_sc_hd__a221o_1
XFILLER_220_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19152_ _19649_/CLK _19152_/D vssd1 vssd1 vccd1 vccd1 _19152_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16364_ _17663_/A0 _18975_/Q _16385_/S vssd1 vssd1 vccd1 vccd1 _18975_/D sky130_fd_sc_hd__mux2_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ _13576_/A vssd1 vssd1 vccd1 vccd1 _13576_/Y sky130_fd_sc_hd__inv_2
X_10788_ _10785_/X _10787_/X _10399_/A vssd1 vssd1 vccd1 vccd1 _10788_/Y sky130_fd_sc_hd__a21oi_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _18734_/CLK _18103_/D vssd1 vssd1 vccd1 vccd1 _18103_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_185_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15315_ _18571_/Q _15314_/C _18572_/Q vssd1 vssd1 vccd1 vccd1 _15315_/Y sky130_fd_sc_hd__a21oi_1
X_12527_ _12521_/X _12522_/Y _12525_/X _12526_/X vssd1 vssd1 vccd1 vccd1 _12527_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19083_ _19197_/CLK _19083_/D vssd1 vssd1 vccd1 vccd1 _19083_/Q sky130_fd_sc_hd__dfxtp_1
X_16295_ _17693_/A0 _18908_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _18908_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18034_ _19636_/CLK _18034_/D vssd1 vssd1 vccd1 vccd1 _18034_/Q sky130_fd_sc_hd__dfxtp_1
X_15246_ _18569_/Q _15270_/C _15223_/A vssd1 vssd1 vccd1 vccd1 _15247_/B sky130_fd_sc_hd__o21ai_1
X_12458_ _14669_/B _16819_/C vssd1 vssd1 vccd1 vccd1 _12458_/Y sky130_fd_sc_hd__nor2_1
X_11409_ _09089_/Y _11398_/X _11406_/X _11408_/X vssd1 vssd1 vccd1 vccd1 _11409_/Y
+ sky130_fd_sc_hd__o31ai_4
X_12389_ _12389_/A1 _12430_/A _12388_/Y _14001_/C1 vssd1 vssd1 vccd1 vccd1 _17904_/D
+ sky130_fd_sc_hd__o211a_1
X_15177_ _15177_/A _15177_/B vssd1 vssd1 vccd1 vccd1 _15179_/B sky130_fd_sc_hd__xnor2_2
XFILLER_99_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14128_ _17711_/A0 _18067_/Q _14140_/S vssd1 vssd1 vccd1 vccd1 _18067_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18936_ _19647_/CLK _18936_/D vssd1 vssd1 vccd1 vccd1 _18936_/Q sky130_fd_sc_hd__dfxtp_1
X_14059_ _16609_/A0 _18001_/Q _14073_/S vssd1 vssd1 vccd1 vccd1 _18001_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18867_ _19219_/CLK _18867_/D vssd1 vssd1 vccd1 vccd1 _18867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_255_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17818_ _19490_/CLK _17818_/D vssd1 vssd1 vccd1 vccd1 _17818_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_283_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18798_ _19632_/CLK _18798_/D vssd1 vssd1 vccd1 vccd1 _18798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17749_ _18649_/Q vssd1 vssd1 vccd1 vccd1 _18649_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_282_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19419_ _19484_/CLK _19419_/D vssd1 vssd1 vccd1 vccd1 _19419_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_189_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09103_ _08948_/A _08948_/B _09102_/X vssd1 vssd1 vccd1 vccd1 _09103_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_248_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09034_ _09048_/A _09034_/B vssd1 vssd1 vccd1 vccd1 _09326_/A sky130_fd_sc_hd__nor2_4
XFILLER_136_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout800 _16293_/Y vssd1 vssd1 vccd1 vccd1 _16325_/S sky130_fd_sc_hd__buf_12
XFILLER_277_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout811 _14483_/S vssd1 vssd1 vccd1 vccd1 _14485_/S sky130_fd_sc_hd__buf_12
Xfanout1809 _17376_/A vssd1 vssd1 vccd1 vccd1 _14442_/B sky130_fd_sc_hd__clkbuf_4
Xfanout822 _14301_/S vssd1 vssd1 vccd1 vccd1 _14304_/S sky130_fd_sc_hd__buf_12
X_09936_ _19619_/Q _18908_/Q _09937_/S vssd1 vssd1 vccd1 vccd1 _09936_/X sky130_fd_sc_hd__mux2_1
Xfanout833 _11144_/X vssd1 vssd1 vccd1 vccd1 _16476_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout844 _16545_/A0 vssd1 vssd1 vccd1 vccd1 _17711_/A0 sky130_fd_sc_hd__buf_4
XFILLER_113_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout855 _10713_/A2 vssd1 vssd1 vccd1 vccd1 _17714_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_246_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout866 _10341_/A2 vssd1 vssd1 vccd1 vccd1 _16553_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout877 _15832_/A1 vssd1 vssd1 vccd1 vccd1 _16622_/A0 sky130_fd_sc_hd__clkbuf_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09867_ _18845_/Q _18877_/Q _19037_/Q _19005_/Q _09885_/S _17905_/Q vssd1 vssd1 vccd1
+ vccd1 _09867_/X sky130_fd_sc_hd__mux4_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout888 _09984_/A vssd1 vssd1 vccd1 vccd1 _12935_/S sky130_fd_sc_hd__buf_4
XFILLER_258_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout899 _09334_/X vssd1 vssd1 vccd1 vccd1 _17667_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_246_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08818_ _19462_/Q vssd1 vssd1 vccd1 vccd1 _08818_/Y sky130_fd_sc_hd__inv_2
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09798_ _18535_/Q _18410_/Q _09801_/S vssd1 vssd1 vccd1 vccd1 _09798_/X sky130_fd_sc_hd__mux2_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _17802_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _17913_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_226 _18385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _18394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_248 _18731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11760_ _18578_/Q _14349_/B _11770_/B1 _13476_/B vssd1 vssd1 vccd1 vccd1 _11760_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_259 input216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10711_ _12320_/A _10689_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _10711_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11691_ _18268_/Q _11695_/B _11691_/B1 vssd1 vssd1 vccd1 vccd1 _11691_/X sky130_fd_sc_hd__a21o_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10642_ _18555_/Q _18430_/Q _10645_/S vssd1 vssd1 vccd1 vccd1 _10642_/X sky130_fd_sc_hd__mux2_1
X_13430_ _19407_/Q _13654_/A2 _13654_/B1 vssd1 vssd1 vccd1 vccd1 _13430_/X sky130_fd_sc_hd__a21o_1
XFILLER_195_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13361_ _13323_/X _13348_/X _13360_/X _13968_/B2 vssd1 vssd1 vccd1 vccd1 _13361_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10573_ _19123_/Q _19155_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _10573_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15100_ _19391_/Q _15092_/B input177/X _15085_/X _15099_/X vssd1 vssd1 vccd1 vccd1
+ _15101_/D sky130_fd_sc_hd__a311o_1
XFILLER_181_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12312_ _15082_/C _12312_/B vssd1 vssd1 vccd1 vccd1 _12312_/X sky130_fd_sc_hd__or2_4
X_16080_ _16096_/A1 _16079_/Y _17725_/C1 vssd1 vssd1 vccd1 vccd1 _18742_/D sky130_fd_sc_hd__a21oi_1
XFILLER_177_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13292_ _08892_/X _13292_/A2 _13291_/X _12762_/B _17931_/Q vssd1 vssd1 vccd1 vccd1
+ _13293_/B sky130_fd_sc_hd__a32o_1
XFILLER_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15031_ _18520_/Q input197/X _15038_/S vssd1 vssd1 vccd1 vccd1 _18520_/D sky130_fd_sc_hd__mux2_1
X_12243_ _12243_/A _12248_/C vssd1 vssd1 vccd1 vccd1 _12243_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12174_ _17854_/Q _12176_/C _12173_/Y vssd1 vssd1 vccd1 vccd1 _17854_/D sky130_fd_sc_hd__o21a_1
XFILLER_218_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11125_ _11352_/A1 _19603_/Q _19571_/Q _11125_/B2 vssd1 vssd1 vccd1 vccd1 _11125_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16982_ _17555_/B _17591_/C _17381_/B vssd1 vssd1 vccd1 vccd1 _17003_/B sky130_fd_sc_hd__nor3_4
X_18721_ _18772_/CLK _18721_/D vssd1 vssd1 vccd1 vccd1 _18721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15933_ _18686_/Q _15948_/A2 _15923_/C _15932_/X _15945_/C1 vssd1 vssd1 vccd1 vccd1
+ _15933_/X sky130_fd_sc_hd__a221o_1
XFILLER_249_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ _13515_/A vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__inv_2
XFILLER_114_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10007_ _11567_/S _10006_/X _10005_/X _11084_/S vssd1 vssd1 vccd1 vccd1 _10007_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_265_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18652_ _18666_/CLK _18652_/D vssd1 vssd1 vccd1 vccd1 _18652_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _18663_/Q _15853_/Y _15906_/B1 vssd1 vssd1 vccd1 vccd1 _15864_/X sky130_fd_sc_hd__a21o_1
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _15086_/X _17592_/X _17603_/B1 vssd1 vssd1 vccd1 vccd1 _17603_/X sky130_fd_sc_hd__a21o_1
XFILLER_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _14815_/A vssd1 vssd1 vccd1 vccd1 _14815_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_18_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ _19485_/CLK _18583_/D vssd1 vssd1 vccd1 vccd1 _18583_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _15778_/B _15780_/B _15776_/X vssd1 vssd1 vccd1 vccd1 _15796_/B sky130_fd_sc_hd__a21oi_1
XFILLER_251_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _18129_/Q _17539_/C1 _17214_/A _17205_/B _17390_/Y vssd1 vssd1 vccd1 vccd1
+ _17534_/X sky130_fd_sc_hd__a221o_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14746_ input98/X input73/X _14784_/S vssd1 vssd1 vccd1 vccd1 _14746_/X sky130_fd_sc_hd__mux2_8
XFILLER_205_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11958_ _11666_/A _11780_/X _11663_/A vssd1 vssd1 vccd1 vccd1 _14345_/C sky130_fd_sc_hd__a21o_1
XFILLER_251_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10909_ _13600_/S _10909_/B vssd1 vssd1 vccd1 vccd1 _13597_/A sky130_fd_sc_hd__nor2_8
X_17465_ _13443_/B _17475_/A2 _17475_/B1 _17805_/Q _17550_/A vssd1 vssd1 vccd1 vccd1
+ _17465_/X sky130_fd_sc_hd__a221o_1
XFILLER_199_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14677_ _14681_/C _14679_/B _14681_/B _14679_/D vssd1 vssd1 vccd1 vccd1 _14677_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_149_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11889_ _11815_/Y _11875_/Y _11888_/X vssd1 vssd1 vccd1 vccd1 _11890_/C sky130_fd_sc_hd__o21ai_4
X_19204_ _19208_/CLK _19204_/D vssd1 vssd1 vccd1 vccd1 _19204_/Q sky130_fd_sc_hd__dfxtp_1
X_16416_ _16614_/A0 _19025_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _19025_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13628_ _19543_/Q _13921_/S vssd1 vssd1 vccd1 vccd1 _13628_/X sky130_fd_sc_hd__or2_1
X_17396_ _11826_/A _17445_/A2 _17445_/B1 _17791_/Q vssd1 vssd1 vccd1 vccd1 _17396_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_220_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19135_ _19201_/CLK _19135_/D vssd1 vssd1 vccd1 vccd1 _19135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16347_ _18959_/Q _17679_/A0 _16358_/S vssd1 vssd1 vccd1 vccd1 _18959_/D sky130_fd_sc_hd__mux2_1
X_13559_ _19315_/Q _13174_/A _13722_/B1 _13552_/X _13558_/X vssd1 vssd1 vccd1 vccd1
+ _13559_/Y sky130_fd_sc_hd__a2111oi_2
XFILLER_285_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19066_ _19618_/CLK _19066_/D vssd1 vssd1 vccd1 vccd1 _19066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16278_ _17676_/A0 _18892_/Q _16278_/S vssd1 vssd1 vccd1 vccd1 _18892_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18017_ _19587_/CLK _18017_/D vssd1 vssd1 vccd1 vccd1 _18017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput403 _11925_/X vssd1 vssd1 vccd1 vccd1 din0[5] sky130_fd_sc_hd__buf_4
X_15229_ _19462_/Q _19396_/Q vssd1 vssd1 vccd1 vccd1 _15230_/B sky130_fd_sc_hd__nand2_2
Xoutput414 _18484_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[13] sky130_fd_sc_hd__buf_4
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput425 _18494_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[23] sky130_fd_sc_hd__buf_4
XFILLER_173_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput436 _18475_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[4] sky130_fd_sc_hd__buf_4
Xoutput447 _18735_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[2] sky130_fd_sc_hd__buf_4
XFILLER_126_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput458 _18118_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[17] sky130_fd_sc_hd__buf_4
Xoutput469 _18128_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[27] sky130_fd_sc_hd__buf_4
XFILLER_259_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09721_ _18630_/Q _18052_/Q _09724_/S vssd1 vssd1 vccd1 vccd1 _09721_/X sky130_fd_sc_hd__mux2_1
X_18919_ _19630_/CLK _18919_/D vssd1 vssd1 vccd1 vccd1 _18919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09652_ _09652_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09653_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09583_ _10366_/A1 _18138_/Q _18784_/Q _10362_/S _12766_/A0 vssd1 vssd1 vccd1 vccd1
+ _09583_/X sky130_fd_sc_hd__a221o_1
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09017_ _09031_/S _09006_/X _09016_/X vssd1 vssd1 vccd1 vccd1 _09017_/X sky130_fd_sc_hd__a21o_1
XFILLER_152_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1606 _15104_/X vssd1 vssd1 vccd1 vccd1 _17445_/C1 sky130_fd_sc_hd__buf_2
Xfanout1617 _09013_/Y vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_132_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout630 _16843_/X vssd1 vssd1 vccd1 vccd1 _16963_/S sky130_fd_sc_hd__clkbuf_4
Xfanout1628 _08986_/Y vssd1 vssd1 vccd1 vccd1 _09650_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1639 _09012_/A vssd1 vssd1 vccd1 vccd1 _09908_/A1 sky130_fd_sc_hd__buf_4
Xfanout641 _17337_/S vssd1 vssd1 vccd1 vccd1 _17345_/S sky130_fd_sc_hd__buf_4
X_09919_ _09935_/A _09917_/X _09918_/X _09919_/C1 vssd1 vssd1 vccd1 vccd1 _09919_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout652 _17009_/B vssd1 vssd1 vccd1 vccd1 _17043_/B sky130_fd_sc_hd__buf_4
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout663 _12562_/X vssd1 vssd1 vccd1 vccd1 _13064_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_59_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout674 _14996_/A1 vssd1 vssd1 vccd1 vccd1 _15006_/A1 sky130_fd_sc_hd__buf_8
XFILLER_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout685 _13655_/A2 vssd1 vssd1 vccd1 vccd1 _13949_/A2 sky130_fd_sc_hd__buf_4
XFILLER_219_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout696 _12556_/Y vssd1 vssd1 vccd1 vccd1 _13246_/A2 sky130_fd_sc_hd__buf_6
X_12930_ _12810_/A _12812_/X _12935_/S vssd1 vssd1 vccd1 vccd1 _12930_/X sky130_fd_sc_hd__mux2_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12860_/X _15863_/A _12918_/S vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__mux2_1
XFILLER_246_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _16526_/A0 _18407_/Q _14622_/S vssd1 vssd1 vccd1 vccd1 _18407_/D sky130_fd_sc_hd__mux2_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11812_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11812_/X sky130_fd_sc_hd__or2_4
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15580_ _15580_/A _15580_/B _15638_/B vssd1 vssd1 vccd1 vccd1 _15580_/X sky130_fd_sc_hd__or3_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _13462_/A _12784_/Y _12785_/X _12791_/X vssd1 vssd1 vccd1 vccd1 _12792_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_233_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _18374_/Q _14559_/A2 _14559_/B1 input21/X vssd1 vssd1 vccd1 vccd1 _14532_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11743_/A _13083_/A vssd1 vssd1 vccd1 vccd1 _13081_/A sky130_fd_sc_hd__xnor2_4
XFILLER_187_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _17443_/A _17250_/B vssd1 vssd1 vccd1 vccd1 _17250_/Y sky130_fd_sc_hd__nor2_1
X_14462_ _18314_/Q _17666_/A0 _14483_/S vssd1 vssd1 vccd1 vccd1 _18314_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11674_ _11674_/A _13568_/A vssd1 vssd1 vccd1 vccd1 _13566_/A sky130_fd_sc_hd__xor2_4
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16201_ _17698_/A0 _18817_/Q _16222_/S vssd1 vssd1 vccd1 vccd1 _18817_/D sky130_fd_sc_hd__mux2_1
X_13413_ _13390_/S _12738_/Y _13413_/B1 vssd1 vssd1 vccd1 vccd1 _13413_/X sky130_fd_sc_hd__a21o_1
XFILLER_169_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17181_ _17208_/A _17181_/B vssd1 vssd1 vccd1 vccd1 _17493_/A sky130_fd_sc_hd__nand2_1
X_10625_ _10625_/A1 _19577_/Q _09108_/B _19609_/Q vssd1 vssd1 vccd1 vccd1 _10625_/X
+ sky130_fd_sc_hd__o22a_1
X_14393_ _17700_/A0 _18244_/Q _14415_/S vssd1 vssd1 vccd1 vccd1 _18244_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16132_ _16142_/A1 _16131_/Y _16142_/B1 vssd1 vssd1 vccd1 vccd1 _18768_/D sky130_fd_sc_hd__a21oi_1
XFILLER_128_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13344_ _17836_/Q _13821_/B _13343_/X vssd1 vssd1 vccd1 vccd1 _13344_/X sky130_fd_sc_hd__o21a_1
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10556_ _10850_/A1 _19155_/Q _09108_/B _19123_/Q vssd1 vssd1 vccd1 vccd1 _10556_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16063_ _16063_/A _16063_/B _16063_/C vssd1 vssd1 vccd1 vccd1 _16063_/Y sky130_fd_sc_hd__nand3_1
X_13275_ _17834_/Q _13942_/A2 _13942_/B1 _17866_/Q vssd1 vssd1 vccd1 vccd1 _13275_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ _10623_/A _10486_/Y _10473_/Y _10532_/A vssd1 vssd1 vccd1 vccd1 _10487_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_185_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15014_ _17159_/A _15014_/B _15014_/C vssd1 vssd1 vccd1 vccd1 _15014_/Y sky130_fd_sc_hd__nor3_1
X_12226_ _17874_/Q _12226_/B vssd1 vssd1 vccd1 vccd1 _12232_/C sky130_fd_sc_hd__and2_2
XFILLER_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12157_ _17848_/Q _12160_/C _12243_/A vssd1 vssd1 vccd1 vccd1 _12157_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_151_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11108_ _11352_/A1 _18611_/Q _18182_/Q _11353_/B2 vssd1 vssd1 vccd1 vccd1 _11108_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_256_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16965_ _18772_/Q _16965_/A2 _16965_/B1 input238/X _16965_/C1 vssd1 vssd1 vccd1 vccd1
+ _16965_/X sky130_fd_sc_hd__a221o_1
X_12088_ _17919_/Q _12088_/A2 _12087_/X _17328_/A vssd1 vssd1 vccd1 vccd1 _17821_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15916_ _18681_/Q _15943_/A2 _15915_/X _15946_/C1 vssd1 vssd1 vccd1 vccd1 _18681_/D
+ sky130_fd_sc_hd__o211a_1
X_11039_ _11039_/A _11039_/B vssd1 vssd1 vccd1 vccd1 _11039_/Y sky130_fd_sc_hd__nor2_1
X_18704_ _19306_/CLK _18704_/D vssd1 vssd1 vccd1 vccd1 _18704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16896_ _16904_/A _16896_/B vssd1 vssd1 vccd1 vccd1 _19308_/D sky130_fd_sc_hd__and2_1
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18635_ _19076_/CLK _18635_/D vssd1 vssd1 vccd1 vccd1 _18635_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_92_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _16041_/A _16063_/A vssd1 vssd1 vccd1 vccd1 _15853_/B sky130_fd_sc_hd__nor2_8
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18566_ _19525_/CLK _18566_/D vssd1 vssd1 vccd1 vccd1 _18566_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _15776_/X _15778_/B vssd1 vssd1 vccd1 vccd1 _15780_/A sky130_fd_sc_hd__nand2b_1
XFILLER_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17517_ _17517_/A _17517_/B vssd1 vssd1 vccd1 vccd1 _17517_/Y sky130_fd_sc_hd__nand2_1
XFILLER_206_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14729_ _14718_/A _14728_/X _14846_/B1 vssd1 vssd1 vccd1 vccd1 _14729_/Y sky130_fd_sc_hd__o21bai_4
X_18497_ _18501_/CLK _18497_/D vssd1 vssd1 vccd1 vccd1 _18497_/Q sky130_fd_sc_hd__dfxtp_1
X_17448_ _17448_/A _17453_/B vssd1 vssd1 vccd1 vccd1 _17448_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17379_ _19487_/Q _17214_/B _17379_/S vssd1 vssd1 vccd1 vccd1 _17380_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19621_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19118_ _19118_/CLK _19118_/D vssd1 vssd1 vccd1 vccd1 _19118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19049_ _19216_/CLK _19049_/D vssd1 vssd1 vccd1 vccd1 _19049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput288 _11963_/X vssd1 vssd1 vccd1 vccd1 addr0[3] sky130_fd_sc_hd__buf_4
Xoutput299 _11915_/X vssd1 vssd1 vccd1 vccd1 addr1[5] sky130_fd_sc_hd__buf_4
XFILLER_88_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09704_ _19039_/Q _19007_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09704_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09635_ _09690_/A _09626_/Y _09630_/Y _08843_/A vssd1 vssd1 vccd1 vccd1 _09635_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_28_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09566_ _09652_/A _09566_/B vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__nor2_1
XFILLER_270_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09497_ _18242_/Q _18817_/Q _09498_/S vssd1 vssd1 vccd1 vccd1 _09497_/X sky130_fd_sc_hd__mux2_1
XFILLER_208_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10410_ _18652_/Q _18074_/Q _19093_/Q _18997_/Q _11379_/S _09136_/S vssd1 vssd1 vccd1
+ vccd1 _10410_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11390_ _09129_/S _11388_/X _11389_/X _11466_/B1 vssd1 vssd1 vccd1 vccd1 _11390_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ _09611_/A _10341_/A2 _10340_/Y _11257_/C1 vssd1 vssd1 vccd1 vccd1 _10342_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_137_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ _15908_/A _12536_/Y _12505_/Y vssd1 vssd1 vccd1 vccd1 _13060_/X sky130_fd_sc_hd__a21o_1
XFILLER_191_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10272_ _17916_/Q _11337_/B _11489_/B1 _10271_/Y vssd1 vssd1 vccd1 vccd1 _10307_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12011_ _17778_/Q _17679_/A0 _12022_/S vssd1 vssd1 vccd1 vccd1 _17778_/D sky130_fd_sc_hd__mux2_1
XFILLER_279_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1403 _09539_/S vssd1 vssd1 vccd1 vccd1 _09542_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_120_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1414 fanout1415/X vssd1 vssd1 vccd1 vccd1 _10090_/S sky130_fd_sc_hd__buf_6
XFILLER_239_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1425 _11403_/S vssd1 vssd1 vccd1 vccd1 _11379_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1436 _10632_/S vssd1 vssd1 vccd1 vccd1 _10557_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1447 _11559_/S1 vssd1 vssd1 vccd1 vccd1 _11311_/C1 sky130_fd_sc_hd__buf_6
Xfanout1458 _09000_/Y vssd1 vssd1 vccd1 vccd1 _09027_/A sky130_fd_sc_hd__buf_4
XFILLER_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1469 fanout1525/X vssd1 vssd1 vccd1 vccd1 fanout1469/X sky130_fd_sc_hd__clkbuf_8
X_16750_ _19269_/Q _16751_/C _19270_/Q vssd1 vssd1 vccd1 vccd1 _16752_/B sky130_fd_sc_hd__a21oi_1
XFILLER_87_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout493 _14667_/X vssd1 vssd1 vccd1 vccd1 _15011_/A2 sky130_fd_sc_hd__buf_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13962_ _13962_/A _13962_/B vssd1 vssd1 vccd1 vccd1 _13962_/Y sky130_fd_sc_hd__nor2_1
XFILLER_246_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15701_ _18128_/Q _15133_/Y _15700_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _15702_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_47_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_79_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19196_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_206_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12913_ _19459_/Q _12529_/Y _12578_/Y _19331_/Q _12912_/X vssd1 vssd1 vccd1 vccd1
+ _12913_/X sky130_fd_sc_hd__a221o_1
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16681_ _19245_/Q _19244_/Q _19241_/Q _19236_/Q vssd1 vssd1 vccd1 vccd1 _16683_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_207_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13893_ _13904_/B _13958_/B _13892_/Y vssd1 vssd1 vccd1 vccd1 _13893_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18420_ _19599_/CLK _18420_/D vssd1 vssd1 vccd1 vccd1 _18420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15632_ _19479_/Q _15631_/Y _15781_/S vssd1 vssd1 vccd1 vccd1 _15632_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12844_ _12448_/D _12840_/X _12843_/X _12792_/X vssd1 vssd1 vccd1 vccd1 _12844_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18351_ _19629_/CLK _18351_/D vssd1 vssd1 vccd1 vccd1 _18351_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15623_/A _15561_/X _15562_/Y _15793_/A2 vssd1 vssd1 vccd1 vccd1 _15563_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12775_ _19457_/Q _12529_/Y _12578_/Y _19329_/Q _12774_/X vssd1 vssd1 vccd1 vccd1
+ _12775_/X sky130_fd_sc_hd__a221o_1
XFILLER_15_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17302_ _18128_/Q _15717_/B2 _17202_/Y _17289_/B vssd1 vssd1 vccd1 vccd1 _17302_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14514_ _17716_/A0 _18364_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _18364_/D sky130_fd_sc_hd__mux2_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11726_ _18778_/Q _11726_/B vssd1 vssd1 vccd1 vccd1 _11726_/X sky130_fd_sc_hd__and2_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _18778_/CLK _18282_/D vssd1 vssd1 vccd1 vccd1 _18282_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _19473_/Q _19407_/Q vssd1 vssd1 vccd1 vccd1 _15496_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17233_ _18105_/Q _17382_/A _17413_/A _17241_/B vssd1 vssd1 vccd1 vccd1 _17233_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14445_ _18584_/Q _14449_/B vssd1 vssd1 vccd1 vccd1 _18297_/D sky130_fd_sc_hd__and2_1
XFILLER_30_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11657_ _12264_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _12837_/B sky130_fd_sc_hd__nand2_8
XFILLER_128_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10608_ _10606_/X _10607_/X _08947_/B vssd1 vssd1 vccd1 vccd1 _10608_/X sky130_fd_sc_hd__a21o_1
X_17164_ _19406_/Q fanout534/X _17462_/A _17212_/B2 vssd1 vssd1 vccd1 vccd1 _17165_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14376_ _18228_/Q _10532_/B _14383_/S vssd1 vssd1 vccd1 vccd1 _18228_/D sky130_fd_sc_hd__mux2_1
X_11588_ _11583_/Y _11587_/X _11588_/B1 vssd1 vssd1 vccd1 vccd1 _11588_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16115_ _18760_/Q _16139_/B vssd1 vssd1 vccd1 vccd1 _16115_/Y sky130_fd_sc_hd__nand2_1
X_13327_ _13397_/C _13327_/B vssd1 vssd1 vccd1 vccd1 _13327_/X sky130_fd_sc_hd__or2_1
XFILLER_143_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10539_ _10866_/S _10538_/X _10537_/X vssd1 vssd1 vccd1 vccd1 _10539_/Y sky130_fd_sc_hd__o21ai_1
X_17095_ _19381_/Q _17107_/B vssd1 vssd1 vccd1 vccd1 _17095_/X sky130_fd_sc_hd__or2_1
XFILLER_171_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16046_ _16046_/A _16046_/B vssd1 vssd1 vccd1 vccd1 _18734_/D sky130_fd_sc_hd__and2_1
XFILLER_143_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13258_ _13258_/A _13312_/A vssd1 vssd1 vccd1 vccd1 _13258_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12209_ _16811_/A _12209_/B _12210_/B vssd1 vssd1 vccd1 vccd1 _17867_/D sky130_fd_sc_hd__nor3_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13189_ _13225_/C _13189_/B vssd1 vssd1 vccd1 vccd1 _14143_/C sky130_fd_sc_hd__nor2_1
XFILLER_285_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17997_ _19599_/CLK _17997_/D vssd1 vssd1 vccd1 vccd1 _17997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16948_ _16960_/A _16948_/B vssd1 vssd1 vccd1 vccd1 _19321_/D sky130_fd_sc_hd__and2_1
XFILLER_38_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16879_ _19304_/Q _17575_/A _16967_/S vssd1 vssd1 vccd1 vccd1 _16880_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09420_ _10366_/A1 _18946_/Q _18211_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09420_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18618_ _19641_/CLK _18618_/D vssd1 vssd1 vccd1 vccd1 _18618_/Q sky130_fd_sc_hd__dfxtp_1
X_19598_ _19612_/CLK _19598_/D vssd1 vssd1 vccd1 vccd1 _19598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_252_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09351_ _18244_/Q _18819_/Q _18447_/Q _18348_/Q _10099_/S _08843_/A vssd1 vssd1 vccd1
+ vccd1 _09351_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18549_ _19148_/CLK _18549_/D vssd1 vssd1 vccd1 vccd1 _18549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09282_ _18852_/Q _18884_/Q _09306_/S vssd1 vssd1 vccd1 vccd1 _09282_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08997_ _09043_/A _11556_/B _09245_/C vssd1 vssd1 vccd1 vccd1 _08997_/X sky130_fd_sc_hd__or3_1
XFILLER_272_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09618_ _10323_/A1 _18209_/Q _09688_/S _18944_/Q vssd1 vssd1 vccd1 vccd1 _09618_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_284_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ _10888_/X _10889_/X _11361_/S vssd1 vssd1 vccd1 vccd1 _10890_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09549_ _09553_/A _09540_/Y _09544_/Y _15129_/B2 vssd1 vssd1 vccd1 vccd1 _09549_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_93_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12560_ _12560_/A _12560_/B vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _11511_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11511_/Y sky130_fd_sc_hd__nand2_1
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_197_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19649_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12491_ _12491_/A _12572_/A _12553_/C vssd1 vssd1 vccd1 vccd1 _12548_/A sky130_fd_sc_hd__or3_4
XFILLER_196_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14230_ _18113_/Q _14260_/B vssd1 vssd1 vccd1 vccd1 _14230_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_126_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19320_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11442_ _09141_/A _15380_/A _11441_/X vssd1 vssd1 vccd1 vccd1 _12597_/B sky130_fd_sc_hd__o21ai_4
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11373_ _09050_/X _09574_/B _11372_/Y _09030_/X vssd1 vssd1 vccd1 vccd1 _11373_/X
+ sky130_fd_sc_hd__o22a_1
X_14161_ _18740_/Q _16054_/A _16034_/S _18741_/Q vssd1 vssd1 vccd1 vccd1 _14164_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10324_ _10322_/X _10323_/X _11173_/S vssd1 vssd1 vccd1 vccd1 _10324_/X sky130_fd_sc_hd__mux2_1
X_13112_ _19367_/Q _13247_/A2 _13110_/X _13111_/X _13247_/C1 vssd1 vssd1 vccd1 vccd1
+ _13112_/X sky130_fd_sc_hd__o221a_4
X_14092_ _17708_/A0 _18032_/Q _14098_/S vssd1 vssd1 vccd1 vccd1 _18032_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10255_ _10243_/A _10250_/X _10252_/X _10254_/X _09264_/S vssd1 vssd1 vccd1 vccd1
+ _10255_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_140_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17920_ _19650_/CLK _17920_/D vssd1 vssd1 vccd1 vccd1 _17920_/Q sky130_fd_sc_hd__dfxtp_4
X_13043_ _13136_/S _13042_/X _13040_/X vssd1 vssd1 vccd1 vccd1 _13043_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_285_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1200 _13230_/A1 vssd1 vssd1 vccd1 vccd1 _13316_/B sky130_fd_sc_hd__buf_8
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1211 _14154_/B1 vssd1 vssd1 vccd1 vccd1 _12835_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17851_ _19310_/CLK _17851_/D vssd1 vssd1 vccd1 vccd1 _17851_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_182_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10186_ _10250_/S _10181_/X _10185_/X vssd1 vssd1 vccd1 vccd1 _10186_/X sky130_fd_sc_hd__o21a_1
XFILLER_239_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1222 _13899_/A vssd1 vssd1 vccd1 vccd1 _15452_/A sky130_fd_sc_hd__buf_4
Xfanout1233 _12265_/Y vssd1 vssd1 vccd1 vccd1 _13966_/C1 sky130_fd_sc_hd__clkbuf_8
Xfanout1244 _08944_/Y vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__buf_8
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16802_ _19289_/Q _16802_/B vssd1 vssd1 vccd1 vccd1 _16807_/C sky130_fd_sc_hd__and2_2
Xfanout1255 _10905_/S vssd1 vssd1 vccd1 vccd1 _13545_/A sky130_fd_sc_hd__buf_2
XFILLER_182_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17782_ _19638_/CLK _17782_/D vssd1 vssd1 vccd1 vccd1 _17782_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1266 _09866_/B vssd1 vssd1 vccd1 vccd1 _13185_/A sky130_fd_sc_hd__buf_6
X_14994_ _18131_/Q _14994_/B vssd1 vssd1 vccd1 vccd1 _14994_/X sky130_fd_sc_hd__or2_1
Xfanout1277 _11715_/B vssd1 vssd1 vccd1 vccd1 _14875_/B1 sky130_fd_sc_hd__buf_6
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1288 _15037_/S vssd1 vssd1 vccd1 vccd1 _15024_/S sky130_fd_sc_hd__buf_2
XFILLER_120_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1299 _12786_/X vssd1 vssd1 vccd1 vccd1 _15789_/A1 sky130_fd_sc_hd__buf_6
X_16733_ _19263_/Q _16736_/D _19264_/Q vssd1 vssd1 vccd1 vccd1 _16735_/B sky130_fd_sc_hd__a21oi_1
X_19521_ _19521_/CLK _19521_/D vssd1 vssd1 vccd1 vccd1 _19521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13945_ _17886_/Q _13945_/A2 _13943_/X _13945_/B2 vssd1 vssd1 vccd1 vccd1 _13945_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19452_ _19453_/CLK _19452_/D vssd1 vssd1 vccd1 vccd1 _19452_/Q sky130_fd_sc_hd__dfxtp_1
X_16664_ _19243_/Q _19242_/Q _16664_/C vssd1 vssd1 vccd1 vccd1 _16670_/C sky130_fd_sc_hd__and3_1
XFILLER_234_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13876_ _17852_/Q _13944_/B _12548_/X vssd1 vssd1 vccd1 vccd1 _13876_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18403_ _19464_/CLK _18403_/D vssd1 vssd1 vccd1 vccd1 _18403_/Q sky130_fd_sc_hd__dfxtp_4
X_15615_ _18584_/Q _15800_/A2 _15607_/X _15614_/X _17368_/A vssd1 vssd1 vccd1 vccd1
+ _18584_/D sky130_fd_sc_hd__o221a_1
X_12827_ _12820_/X _12826_/Y _13130_/A vssd1 vssd1 vccd1 vccd1 _12827_/X sky130_fd_sc_hd__mux2_1
X_19383_ _19546_/CLK _19383_/D vssd1 vssd1 vccd1 vccd1 _19383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16595_ _16595_/A0 _19198_/Q _16623_/S vssd1 vssd1 vccd1 vccd1 _19198_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18334_ _19613_/CLK _18334_/D vssd1 vssd1 vccd1 vccd1 _18334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ _15538_/X _15539_/X _15545_/X _15782_/A1 _15633_/C1 vssd1 vssd1 vccd1 vccd1
+ _15546_/X sky130_fd_sc_hd__a221o_1
X_12758_ _11650_/B _13358_/A1 _12756_/Y _10065_/B _12757_/X vssd1 vssd1 vccd1 vccd1
+ _12758_/X sky130_fd_sc_hd__o221a_1
XFILLER_203_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18265_ _19225_/CLK _18265_/D vssd1 vssd1 vccd1 vccd1 _18265_/Q sky130_fd_sc_hd__dfxtp_1
X_11709_ _18518_/Q _11708_/X _11711_/A vssd1 vssd1 vccd1 vccd1 _11715_/A sky130_fd_sc_hd__o21a_1
XFILLER_187_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15477_ _18578_/Q _15447_/B _15469_/Y _15476_/X _17350_/A vssd1 vssd1 vccd1 vccd1
+ _18578_/D sky130_fd_sc_hd__o221a_1
XFILLER_202_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12689_ _09984_/B _12660_/B _13911_/A vssd1 vssd1 vccd1 vccd1 _12689_/X sky130_fd_sc_hd__mux2_1
X_17216_ _19423_/Q _17120_/Y _17215_/X vssd1 vssd1 vccd1 vccd1 _19423_/D sky130_fd_sc_hd__o21ba_1
X_14428_ _18567_/Q _16046_/A vssd1 vssd1 vccd1 vccd1 _18280_/D sky130_fd_sc_hd__and2_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18196_ _19639_/CLK _18196_/D vssd1 vssd1 vccd1 vccd1 _18196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ _17255_/A _17147_/B vssd1 vssd1 vccd1 vccd1 _19400_/D sky130_fd_sc_hd__nor2_1
XFILLER_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14359_ _18211_/Q _09437_/B _14380_/S vssd1 vssd1 vccd1 vccd1 _18211_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17078_ _17583_/A _17114_/A2 _17077_/X _17346_/A vssd1 vssd1 vccd1 vccd1 _19372_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08920_ _14350_/A _14488_/B _14306_/C vssd1 vssd1 vccd1 vccd1 _16525_/A sky130_fd_sc_hd__and3_4
X_16029_ _16020_/Y _16028_/X _16027_/X _16052_/A vssd1 vssd1 vccd1 vccd1 _18728_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08851_ _17900_/Q vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__clkinv_2
XFILLER_85_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09403_ _13154_/S _09403_/B vssd1 vssd1 vccd1 vccd1 _13148_/A sky130_fd_sc_hd__and2_4
XFILLER_213_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09334_ _09333_/Y _09332_/X _08945_/X _17928_/Q vssd1 vssd1 vccd1 vccd1 _09334_/X
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09265_ _18245_/Q _18820_/Q _18448_/Q _18349_/Q _09252_/S _12466_/A0 vssd1 vssd1
+ vccd1 vccd1 _09265_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09196_ _12389_/A1 _09195_/X _09194_/X vssd1 vssd1 vccd1 vccd1 _09196_/X sky130_fd_sc_hd__o21a_1
XFILLER_181_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10040_ _10038_/X _10039_/X _10040_/S vssd1 vssd1 vccd1 vccd1 _10041_/B sky130_fd_sc_hd__mux2_1
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11991_ _17758_/Q _16526_/A0 _12013_/S vssd1 vssd1 vccd1 vccd1 _17758_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13730_ _10603_/A _13912_/A2 _13912_/B1 vssd1 vssd1 vccd1 vccd1 _13730_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10942_ _10940_/X _10941_/X _11327_/S vssd1 vssd1 vccd1 vccd1 _10942_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13661_ _13930_/A1 _13647_/Y _13930_/B1 vssd1 vssd1 vccd1 vccd1 _13661_/X sky130_fd_sc_hd__o21a_1
XFILLER_232_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10873_ _11103_/A _11854_/A vssd1 vssd1 vccd1 vccd1 _10873_/Y sky130_fd_sc_hd__nor2_1
XFILLER_220_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15400_ _19469_/Q _15399_/Y _15400_/S vssd1 vssd1 vccd1 vccd1 _15400_/X sky130_fd_sc_hd__mux2_2
XFILLER_188_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _09475_/B _12612_/B vssd1 vssd1 vccd1 vccd1 _12612_/Y sky130_fd_sc_hd__nand2b_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _17679_/A0 _18991_/Q _16391_/S vssd1 vssd1 vccd1 vccd1 _18991_/D sky130_fd_sc_hd__mux2_1
XFILLER_213_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13592_ _19316_/Q _13754_/A2 _13722_/B1 _13585_/X _13591_/X vssd1 vssd1 vccd1 vccd1
+ _13592_/Y sky130_fd_sc_hd__a2111oi_2
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _10027_/A _15382_/B2 _15328_/X _15330_/Y vssd1 vssd1 vccd1 vccd1 _15336_/B
+ sky130_fd_sc_hd__o22a_1
X_12543_ _12544_/A _13167_/A vssd1 vssd1 vccd1 vccd1 _12543_/X sky130_fd_sc_hd__or2_4
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18050_ _18632_/CLK _18050_/D vssd1 vssd1 vccd1 vccd1 _18050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15262_ _15262_/A _15262_/B vssd1 vssd1 vccd1 vccd1 _15365_/A sky130_fd_sc_hd__xor2_2
X_12474_ _12483_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _12474_/Y sky130_fd_sc_hd__nor2_2
XFILLER_200_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17001_ _19337_/Q _17045_/B vssd1 vssd1 vccd1 vccd1 _17001_/X sky130_fd_sc_hd__or2_1
X_14213_ _18278_/Q _14252_/B _14212_/X _16046_/A vssd1 vssd1 vccd1 vccd1 _18104_/D
+ sky130_fd_sc_hd__o211a_1
X_11425_ _11506_/A1 _18952_/Q _18217_/Q _10426_/S vssd1 vssd1 vccd1 vccd1 _11425_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15193_ _18566_/Q _15351_/A2 _15191_/X _15192_/Y _14430_/B vssd1 vssd1 vccd1 vccd1
+ _18566_/D sky130_fd_sc_hd__o221a_1
XFILLER_165_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_7 _18275_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14144_ _14144_/A _14144_/B _13261_/X _13226_/Y vssd1 vssd1 vccd1 vccd1 _14145_/C
+ sky130_fd_sc_hd__or4bb_1
X_11356_ _11356_/A _11356_/B vssd1 vssd1 vccd1 vccd1 _11356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10307_ _10307_/A _12658_/B vssd1 vssd1 vccd1 vccd1 _10308_/A sky130_fd_sc_hd__and2_2
X_18952_ _19612_/CLK _18952_/D vssd1 vssd1 vccd1 vccd1 _18952_/Q sky130_fd_sc_hd__dfxtp_1
X_14075_ _17658_/A _16426_/A vssd1 vssd1 vccd1 vccd1 _14075_/Y sky130_fd_sc_hd__nand2_8
XFILLER_112_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11287_ _11282_/Y _11286_/Y _08950_/A vssd1 vssd1 vccd1 vccd1 _11287_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_94_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18772_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17903_ _18817_/CLK _17903_/D vssd1 vssd1 vccd1 vccd1 _17903_/Q sky130_fd_sc_hd__dfxtp_2
X_13026_ _13930_/A1 _13008_/Y _13253_/B1 vssd1 vssd1 vccd1 vccd1 _13027_/C sky130_fd_sc_hd__o21ai_1
X_10238_ _17948_/Q _11451_/A2 _10237_/X _11451_/B2 vssd1 vssd1 vccd1 vccd1 _10238_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_105_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18883_ _19203_/CLK _18883_/D vssd1 vssd1 vccd1 vccd1 _18883_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1030 _09662_/X vssd1 vssd1 vccd1 vccd1 _16530_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_267_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1041 _09085_/X vssd1 vssd1 vccd1 vccd1 _11411_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_23_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19195_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10169_ _10167_/X _10168_/X _10169_/S vssd1 vssd1 vccd1 vccd1 _10169_/X sky130_fd_sc_hd__mux2_1
X_17834_ _19327_/CLK _17834_/D vssd1 vssd1 vccd1 vccd1 _17834_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1052 _17603_/B1 vssd1 vssd1 vccd1 vccd1 _17623_/B1 sky130_fd_sc_hd__buf_6
Xfanout1063 _13958_/B vssd1 vssd1 vccd1 vccd1 _13861_/A sky130_fd_sc_hd__buf_2
XFILLER_282_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1074 _14027_/A2 vssd1 vssd1 vccd1 vccd1 _14034_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_66_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1085 _17661_/A0 vssd1 vssd1 vccd1 vccd1 _17694_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_266_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1096 _11624_/A1 vssd1 vssd1 vccd1 vccd1 _11210_/A1 sky130_fd_sc_hd__buf_12
XFILLER_282_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17765_ _19614_/CLK _17765_/D vssd1 vssd1 vccd1 vccd1 _17765_/Q sky130_fd_sc_hd__dfxtp_1
X_14977_ input63/X input99/X _15007_/S vssd1 vssd1 vccd1 vccd1 _14978_/A sky130_fd_sc_hd__mux2_2
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19504_ _19552_/CLK _19504_/D vssd1 vssd1 vccd1 vccd1 _19504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16716_ _16808_/A _16722_/C vssd1 vssd1 vccd1 vccd1 _16716_/Y sky130_fd_sc_hd__nor2_1
X_13928_ _13928_/A1 _13918_/X _13927_/X vssd1 vssd1 vccd1 vccd1 _13928_/X sky130_fd_sc_hd__a21o_4
X_17696_ _17696_/A0 _19622_/Q _17719_/S vssd1 vssd1 vccd1 vccd1 _19622_/D sky130_fd_sc_hd__mux2_1
XFILLER_263_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16647_ _19238_/Q _16649_/C _16780_/B1 vssd1 vssd1 vccd1 vccd1 _16648_/B sky130_fd_sc_hd__o21ai_1
X_19435_ _19466_/CLK _19435_/D vssd1 vssd1 vccd1 vccd1 _19435_/Q sky130_fd_sc_hd__dfxtp_2
X_13859_ _17531_/A _13861_/A vssd1 vssd1 vccd1 vccd1 _13859_/X sky130_fd_sc_hd__or2_1
XFILLER_63_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19366_ _19470_/CLK _19366_/D vssd1 vssd1 vccd1 vccd1 _19366_/Q sky130_fd_sc_hd__dfxtp_1
X_16578_ _16611_/A0 _19182_/Q _16585_/S vssd1 vssd1 vccd1 vccd1 _19182_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18317_ _19126_/CLK _18317_/D vssd1 vssd1 vccd1 vccd1 _18317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15529_ _12320_/B _15452_/A _15484_/A vssd1 vssd1 vccd1 vccd1 _15531_/B sky130_fd_sc_hd__o21a_1
XFILLER_124_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19297_ _19326_/CLK _19297_/D vssd1 vssd1 vccd1 vccd1 _19297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09050_ _11141_/A _09050_/B vssd1 vssd1 vccd1 vccd1 _09050_/X sky130_fd_sc_hd__or2_4
XFILLER_187_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18248_ _19629_/CLK _18248_/D vssd1 vssd1 vccd1 vccd1 _18248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18179_ _19216_/CLK _18179_/D vssd1 vssd1 vccd1 vccd1 _18179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09952_ _18595_/Q _18166_/Q _09952_/S vssd1 vssd1 vccd1 vccd1 _09952_/X sky130_fd_sc_hd__mux2_1
XFILLER_249_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08903_ _08903_/A _10275_/S _10364_/B vssd1 vssd1 vccd1 vccd1 _08904_/C sky130_fd_sc_hd__and3_1
XFILLER_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09883_ _18628_/Q _09883_/B vssd1 vssd1 vccd1 vccd1 _09883_/X sky130_fd_sc_hd__or2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08834_ _18108_/Q vssd1 vssd1 vccd1 vccd1 _14220_/A sky130_fd_sc_hd__clkinv_4
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_408 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_419 _15357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09317_ _12600_/A _09317_/B vssd1 vssd1 vccd1 vccd1 _09318_/B sky130_fd_sc_hd__nand2_2
XFILLER_210_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _09247_/Y _09246_/X _08945_/X _17929_/Q vssd1 vssd1 vccd1 vccd1 _09248_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_182_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ _18636_/Q _09179_/B vssd1 vssd1 vccd1 vccd1 _09179_/X sky130_fd_sc_hd__or2_1
XFILLER_135_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11210_ _11210_/A1 _11144_/X _11209_/X vssd1 vssd1 vccd1 vccd1 _15450_/A sky130_fd_sc_hd__a21o_4
XFILLER_108_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12190_ _17860_/Q _12192_/C _12189_/Y vssd1 vssd1 vccd1 vccd1 _17860_/D sky130_fd_sc_hd__o21a_1
XFILLER_108_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ _11141_/A _11141_/B vssd1 vssd1 vccd1 vccd1 _11141_/Y sky130_fd_sc_hd__nor2_1
XFILLER_268_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11072_ _11565_/A1 _18221_/Q _11094_/S _18956_/Q _11559_/S1 vssd1 vssd1 vccd1 vccd1
+ _11072_/X sky130_fd_sc_hd__o221a_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput100 dout0[61] vssd1 vssd1 vccd1 vccd1 input100/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput111 dout1[13] vssd1 vssd1 vccd1 vccd1 input111/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14900_ _18491_/Q _15011_/A2 _14899_/Y _16795_/A vssd1 vssd1 vccd1 vccd1 _18491_/D
+ sky130_fd_sc_hd__a211o_1
Xinput122 dout1[23] vssd1 vssd1 vccd1 vccd1 input122/X sky130_fd_sc_hd__clkbuf_2
X_10023_ _10009_/X _10022_/X _11332_/B1 vssd1 vssd1 vccd1 vccd1 _10023_/X sky130_fd_sc_hd__a21o_2
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _18669_/Q _15949_/A2 _15879_/X _15904_/C1 vssd1 vssd1 vccd1 vccd1 _18669_/D
+ sky130_fd_sc_hd__o211a_1
Xinput133 dout1[33] vssd1 vssd1 vccd1 vccd1 input133/X sky130_fd_sc_hd__buf_2
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput144 dout1[43] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput155 dout1[53] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__buf_2
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 dout1[63] vssd1 vssd1 vccd1 vccd1 input166/X sky130_fd_sc_hd__buf_2
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ _18115_/Q _14994_/B vssd1 vssd1 vccd1 vccd1 _14831_/X sky130_fd_sc_hd__or2_1
Xinput177 irq[15] vssd1 vssd1 vccd1 vccd1 input177/X sky130_fd_sc_hd__clkbuf_4
XFILLER_248_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 jtag_tdi vssd1 vssd1 vccd1 vccd1 _15854_/A sky130_fd_sc_hd__buf_12
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput199 localMemory_wb_adr_i[18] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__clkbuf_2
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _17550_/A _17550_/B vssd1 vssd1 vccd1 vccd1 _17550_/Y sky130_fd_sc_hd__nor2_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ _18108_/Q _14801_/B _14690_/Y _14761_/X vssd1 vssd1 vccd1 vccd1 _14762_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ _18736_/Q _11973_/X _11972_/X vssd1 vssd1 vccd1 vccd1 _15845_/B sky130_fd_sc_hd__o21a_2
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16501_ _16501_/A0 _19107_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _19107_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13713_ _17847_/Q _13846_/B _12548_/X vssd1 vssd1 vccd1 vccd1 _13713_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _11572_/A1 _19573_/Q _10940_/S _19605_/Q _11311_/C1 vssd1 vssd1 vccd1 vccd1
+ _10925_/X sky130_fd_sc_hd__o221a_1
X_17481_ _18580_/Q _17544_/A _08883_/A vssd1 vssd1 vccd1 vccd1 _17481_/X sky130_fd_sc_hd__o21a_1
X_14693_ _14417_/C _12276_/B _14692_/X vssd1 vssd1 vccd1 vccd1 _14693_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16432_ _19040_/Q _16597_/A0 _16454_/S vssd1 vssd1 vccd1 vccd1 _19040_/D sky130_fd_sc_hd__mux2_1
X_19220_ _19642_/CLK _19220_/D vssd1 vssd1 vccd1 vccd1 _19220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_141_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19231_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13644_ _15133_/A _13640_/X _13643_/X _13869_/B2 vssd1 vssd1 vccd1 vccd1 _13644_/Y
+ sky130_fd_sc_hd__a22oi_4
X_10856_ _10866_/S _19183_/Q _10856_/C vssd1 vssd1 vccd1 vccd1 _10856_/X sky130_fd_sc_hd__and3_1
XFILLER_32_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19151_ _19618_/CLK _19151_/D vssd1 vssd1 vccd1 vccd1 _19151_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16529_/A0 _18974_/Q _16391_/S vssd1 vssd1 vccd1 vccd1 _18974_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13575_ _18120_/Q _13606_/C vssd1 vssd1 vccd1 vccd1 _13576_/A sky130_fd_sc_hd__xnor2_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10930_/S _10786_/X _11570_/B1 vssd1 vssd1 vccd1 vccd1 _10787_/X sky130_fd_sc_hd__o21a_1
X_18102_ _18593_/CLK _18102_/D vssd1 vssd1 vccd1 vccd1 _18102_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _18572_/Q _18571_/Q _15314_/C vssd1 vssd1 vccd1 vccd1 _15342_/B sky130_fd_sc_hd__and3_1
XFILLER_200_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _19392_/Q _12575_/A _12577_/B vssd1 vssd1 vccd1 vccd1 _12526_/X sky130_fd_sc_hd__or3_1
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19082_ _19114_/CLK _19082_/D vssd1 vssd1 vccd1 vccd1 _19082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16294_ _17692_/A0 _18907_/Q _16325_/S vssd1 vssd1 vccd1 vccd1 _18907_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18033_ _19635_/CLK _18033_/D vssd1 vssd1 vccd1 vccd1 _18033_/Q sky130_fd_sc_hd__dfxtp_1
X_15245_ _18569_/Q _15270_/C vssd1 vssd1 vccd1 vccd1 _15271_/B sky130_fd_sc_hd__and2_1
X_12457_ _14681_/C _12457_/B vssd1 vssd1 vccd1 vccd1 _16819_/C sky130_fd_sc_hd__nand2b_2
X_11408_ _11387_/X _11390_/X _11407_/X vssd1 vssd1 vccd1 vccd1 _11408_/X sky130_fd_sc_hd__a21o_2
XFILLER_172_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15176_ _14214_/A _15132_/X _15174_/Y _12318_/A _15177_/A vssd1 vssd1 vccd1 vccd1
+ _15200_/A sky130_fd_sc_hd__o221a_1
X_12388_ _12430_/A _12388_/B vssd1 vssd1 vccd1 vccd1 _12388_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ _17677_/A0 _18066_/Q _14139_/S vssd1 vssd1 vccd1 vccd1 _18066_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11339_ _11360_/A1 _19600_/Q _19568_/Q _11340_/B2 vssd1 vssd1 vccd1 vccd1 _11339_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_259_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18935_ _19646_/CLK _18935_/D vssd1 vssd1 vccd1 vccd1 _18935_/Q sky130_fd_sc_hd__dfxtp_1
X_14058_ _17708_/A0 _18000_/Q _14064_/S vssd1 vssd1 vccd1 vccd1 _18000_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13009_ _17828_/Q _13164_/A2 _13164_/B1 _17860_/Q vssd1 vssd1 vccd1 vccd1 _13009_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18866_ _19641_/CLK _18866_/D vssd1 vssd1 vccd1 vccd1 _18866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17817_ _19492_/CLK _17817_/D vssd1 vssd1 vccd1 vccd1 _17817_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_223_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18797_ _19047_/CLK _18797_/D vssd1 vssd1 vccd1 vccd1 _18797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17748_ _18648_/Q vssd1 vssd1 vccd1 vccd1 _18648_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_36_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17679_ _17679_/A0 _19606_/Q _17690_/S vssd1 vssd1 vccd1 vccd1 _19606_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19418_ _19484_/CLK _19418_/D vssd1 vssd1 vccd1 vccd1 _19418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19349_ _19477_/CLK _19349_/D vssd1 vssd1 vccd1 vccd1 _19349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09102_ _09102_/A _09102_/B _09102_/C _09101_/X vssd1 vssd1 vccd1 vccd1 _09102_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_148_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09033_ _11217_/A _09902_/B _09325_/C vssd1 vssd1 vccd1 vccd1 _09033_/X sky130_fd_sc_hd__and3_1
XFILLER_164_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout801 _16165_/S vssd1 vssd1 vccd1 vccd1 _16193_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_277_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09935_ _09935_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09935_/X sky130_fd_sc_hd__or2_1
Xfanout812 _14454_/Y vssd1 vssd1 vccd1 vccd1 _14483_/S sky130_fd_sc_hd__buf_12
XFILLER_264_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout823 _14277_/S vssd1 vssd1 vccd1 vccd1 _14301_/S sky130_fd_sc_hd__buf_12
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout834 _17676_/A0 vssd1 vssd1 vccd1 vccd1 _17709_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout845 _10913_/X vssd1 vssd1 vccd1 vccd1 _16545_/A0 sky130_fd_sc_hd__buf_4
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout856 _10713_/A2 vssd1 vssd1 vccd1 vccd1 _16614_/A0 sky130_fd_sc_hd__clkbuf_2
Xfanout867 _10341_/A2 vssd1 vssd1 vccd1 vccd1 _17686_/A0 sky130_fd_sc_hd__clkbuf_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _14714_/A _09866_/B vssd1 vssd1 vccd1 vccd1 _09866_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout878 _16490_/A0 vssd1 vssd1 vccd1 vccd1 _17722_/A0 sky130_fd_sc_hd__clkbuf_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout889 _09946_/X vssd1 vssd1 vccd1 vccd1 _09984_/A sky130_fd_sc_hd__buf_8
XFILLER_285_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08817_ _19490_/Q vssd1 vssd1 vccd1 vccd1 _08817_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09797_ _18310_/Q _17761_/Q _09797_/S vssd1 vssd1 vccd1 vccd1 _09797_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_205 _18777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_216 _17913_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_227 _18386_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_238 _18394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 _18506_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10707_/X _10709_/X _10326_/A vssd1 vssd1 vccd1 vccd1 _10710_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _18203_/Q _14525_/A vssd1 vssd1 vccd1 vccd1 _11690_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10641_ _18330_/Q _17781_/Q _10645_/S vssd1 vssd1 vccd1 vccd1 _10641_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13360_ _13349_/Y _13352_/Y _13359_/X _12442_/C vssd1 vssd1 vccd1 vccd1 _13360_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10572_ _18072_/Q _10816_/A2 _10571_/X _10643_/S vssd1 vssd1 vccd1 vccd1 _10572_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12311_ _12311_/A vssd1 vssd1 vccd1 vccd1 _12312_/B sky130_fd_sc_hd__clkinv_2
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13291_ _13421_/A _13258_/A _12448_/D _13270_/X _13290_/X vssd1 vssd1 vccd1 vccd1
+ _13291_/X sky130_fd_sc_hd__a221o_1
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15030_ _18519_/Q input196/X _15037_/S vssd1 vssd1 vccd1 vccd1 _18519_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12242_ _17880_/Q _12242_/B vssd1 vssd1 vccd1 vccd1 _12248_/C sky130_fd_sc_hd__and2_2
XFILLER_181_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12173_ _17854_/Q _12176_/C _12203_/A vssd1 vssd1 vccd1 vccd1 _12173_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_218_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11124_ _18549_/Q _18424_/Q _18033_/Q _18001_/Q _11125_/B2 _11338_/S1 vssd1 vssd1
+ vccd1 vccd1 _11124_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16981_ _16981_/A _16981_/B _16840_/B vssd1 vssd1 vccd1 vccd1 _17381_/B sky130_fd_sc_hd__or3b_4
XFILLER_110_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18720_ _18772_/CLK _18720_/D vssd1 vssd1 vccd1 vccd1 _18720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15932_ input3/X input269/X _15947_/S vssd1 vssd1 vccd1 vccd1 _15932_/X sky130_fd_sc_hd__mux2_1
XFILLER_277_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ _11518_/B2 _16610_/A0 _11054_/X _11055_/B2 vssd1 vssd1 vccd1 vccd1 _13515_/A
+ sky130_fd_sc_hd__o2bb2a_4
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10006_ _18532_/Q _18407_/Q _11147_/S vssd1 vssd1 vccd1 vccd1 _10006_/X sky130_fd_sc_hd__mux2_1
X_15863_ _15863_/A _15905_/B _15905_/C vssd1 vssd1 vccd1 vccd1 _15863_/X sky130_fd_sc_hd__and3_1
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18651_ _19092_/CLK _18651_/D vssd1 vssd1 vccd1 vccd1 _18651_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14814_ input46/X input81/X _14844_/S vssd1 vssd1 vccd1 vccd1 _14815_/A sky130_fd_sc_hd__mux2_2
X_17602_ _19542_/Q _17624_/A2 _17591_/X _17181_/B _17601_/X vssd1 vssd1 vccd1 vccd1
+ _19542_/D sky130_fd_sc_hd__o221a_1
XFILLER_92_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18582_ _19444_/CLK _18582_/D vssd1 vssd1 vccd1 vccd1 _18582_/Q sky130_fd_sc_hd__dfxtp_4
X_15794_ _15789_/X _15792_/X _15793_/Y vssd1 vssd1 vccd1 vccd1 _15794_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _14865_/A1 _14744_/X _14865_/B1 vssd1 vssd1 vccd1 vccd1 _14745_/Y sky130_fd_sc_hd__o21ai_2
X_17533_ _17533_/A _17538_/A vssd1 vssd1 vccd1 vccd1 _17533_/Y sky130_fd_sc_hd__nand2_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11957_ _19229_/Q _11959_/A2 _14344_/C _11959_/B2 vssd1 vssd1 vccd1 vccd1 _11957_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_189_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10908_ _12641_/A _10908_/B vssd1 vssd1 vccd1 vccd1 _10909_/B sky130_fd_sc_hd__nor2_4
XFILLER_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17464_ _19504_/Q _17462_/B _17463_/X _17352_/A vssd1 vssd1 vccd1 vccd1 _19504_/D
+ sky130_fd_sc_hd__o211a_1
X_14676_ _14688_/C vssd1 vssd1 vccd1 vccd1 _14679_/D sky130_fd_sc_hd__inv_2
XFILLER_33_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11888_ _11816_/X _11875_/A _11901_/B _11850_/X vssd1 vssd1 vccd1 vccd1 _11888_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_60_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19203_ _19203_/CLK _19203_/D vssd1 vssd1 vccd1 vccd1 _19203_/Q sky130_fd_sc_hd__dfxtp_1
X_16415_ _16580_/A0 _19024_/Q _16420_/S vssd1 vssd1 vccd1 vccd1 _19024_/D sky130_fd_sc_hd__mux2_1
X_13627_ _17876_/Q _13747_/A2 _13625_/X _13682_/B2 vssd1 vssd1 vccd1 vccd1 _13627_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17395_ _19490_/Q _17423_/B _17393_/X _17394_/Y _17328_/A vssd1 vssd1 vccd1 vccd1
+ _19490_/D sky130_fd_sc_hd__o221a_1
X_10839_ _19087_/Q _10840_/S _10838_/X _10918_/C1 vssd1 vssd1 vccd1 vccd1 _10839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16346_ _18958_/Q _16545_/A0 _16358_/S vssd1 vssd1 vccd1 vccd1 _18958_/D sky130_fd_sc_hd__mux2_1
X_19134_ _19134_/CLK _19134_/D vssd1 vssd1 vccd1 vccd1 _19134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13558_ _19379_/Q _13884_/A2 _13556_/X _13557_/X _13884_/C1 vssd1 vssd1 vccd1 vccd1
+ _13558_/X sky130_fd_sc_hd__o221a_4
XFILLER_121_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19065_ _19647_/CLK _19065_/D vssd1 vssd1 vccd1 vccd1 _19065_/Q sky130_fd_sc_hd__dfxtp_1
X_12509_ _12577_/A _12579_/A vssd1 vssd1 vccd1 vccd1 _12575_/A sky130_fd_sc_hd__or2_4
XFILLER_145_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16277_ _16608_/A0 _18891_/Q _16288_/S vssd1 vssd1 vccd1 vccd1 _18891_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13489_ _12835_/A _13390_/X _13391_/Y _13863_/B2 _13488_/X vssd1 vssd1 vccd1 vccd1
+ _13489_/X sky130_fd_sc_hd__o221a_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18016_ _19197_/CLK _18016_/D vssd1 vssd1 vccd1 vccd1 _18016_/Q sky130_fd_sc_hd__dfxtp_1
X_15228_ _19462_/Q _19396_/Q vssd1 vssd1 vccd1 vccd1 _15228_/Y sky130_fd_sc_hd__nor2_2
XFILLER_126_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput404 _11926_/X vssd1 vssd1 vccd1 vccd1 din0[6] sky130_fd_sc_hd__buf_4
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput415 _18485_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[14] sky130_fd_sc_hd__buf_4
Xoutput426 _18495_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[24] sky130_fd_sc_hd__buf_4
Xoutput437 _18476_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[5] sky130_fd_sc_hd__buf_4
XFILLER_160_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput448 _18736_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[3] sky130_fd_sc_hd__buf_4
XFILLER_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15159_ _15149_/Y _15156_/X _15307_/B vssd1 vssd1 vccd1 vccd1 _15159_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput459 _18119_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[18] sky130_fd_sc_hd__buf_4
XFILLER_102_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09720_ _18020_/Q _17988_/Q _09720_/S vssd1 vssd1 vccd1 vccd1 _09720_/X sky130_fd_sc_hd__mux2_1
X_18918_ _19629_/CLK _18918_/D vssd1 vssd1 vccd1 vccd1 _18918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09651_ input110/X input145/X _09651_/S vssd1 vssd1 vccd1 vccd1 _09652_/B sky130_fd_sc_hd__mux2_4
XFILLER_283_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18849_ _18881_/CLK _18849_/D vssd1 vssd1 vccd1 vccd1 _18849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09582_ _18848_/Q _18880_/Q _10362_/S vssd1 vssd1 vccd1 vccd1 _09582_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09016_ _09027_/A _09009_/X _09012_/X _09015_/X vssd1 vssd1 vccd1 vccd1 _09016_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1607 _17527_/A1 vssd1 vssd1 vccd1 vccd1 _17544_/A sky130_fd_sc_hd__buf_4
XFILLER_278_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1618 _09013_/Y vssd1 vssd1 vccd1 vccd1 _09574_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout620 _17158_/B2 vssd1 vssd1 vccd1 vccd1 _17212_/B2 sky130_fd_sc_hd__buf_6
Xfanout631 _12744_/Y vssd1 vssd1 vccd1 vccd1 _13197_/B1 sky130_fd_sc_hd__buf_4
Xfanout1629 _12024_/A vssd1 vssd1 vccd1 vccd1 _12442_/B sky130_fd_sc_hd__buf_12
XFILLER_132_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09918_ _09457_/B _19068_/Q _18972_/Q _11167_/B _10337_/S1 vssd1 vssd1 vccd1 vccd1
+ _09918_/X sky130_fd_sc_hd__o221a_1
Xfanout642 _17108_/A2 vssd1 vssd1 vccd1 vccd1 _17116_/A2 sky130_fd_sc_hd__buf_6
Xfanout653 _17003_/B vssd1 vssd1 vccd1 vccd1 _17009_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_265_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout664 _13654_/A2 vssd1 vssd1 vccd1 vccd1 _13948_/A2 sky130_fd_sc_hd__buf_4
XFILLER_219_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout675 _14694_/X vssd1 vssd1 vccd1 vccd1 _14996_/A1 sky130_fd_sc_hd__buf_4
XFILLER_258_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout686 _12560_/B vssd1 vssd1 vccd1 vccd1 _13655_/A2 sky130_fd_sc_hd__buf_4
XFILLER_246_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout697 _12545_/Y vssd1 vssd1 vccd1 vccd1 _13943_/B1 sky130_fd_sc_hd__buf_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09849_ _09857_/A1 _09845_/X _09848_/X _09106_/B vssd1 vssd1 vccd1 vccd1 _09849_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ input272/X _12575_/Y _12859_/X vssd1 vssd1 vccd1 vccd1 _12860_/X sky130_fd_sc_hd__a21o_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11859_/A _11846_/B vssd1 vssd1 vccd1 vccd1 _11811_/Y sky130_fd_sc_hd__nor2_2
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _13421_/A _11826_/A _12761_/B _12790_/Y _13185_/A vssd1 vssd1 vccd1 vccd1
+ _12791_/X sky130_fd_sc_hd__a221o_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14576_/A _14530_/B vssd1 vssd1 vccd1 vccd1 _18373_/D sky130_fd_sc_hd__or2_1
XFILLER_242_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _09560_/X _11742_/B vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__and2b_4
XFILLER_202_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _18313_/Q _17665_/A0 _14483_/S vssd1 vssd1 vccd1 vccd1 _18313_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11673_ _11673_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _13568_/A sky130_fd_sc_hd__and2_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16200_ _17697_/A0 _18816_/Q _16222_/S vssd1 vssd1 vccd1 vccd1 _18816_/D sky130_fd_sc_hd__mux2_1
XFILLER_169_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13412_ _13958_/B _14147_/A _13892_/B1 vssd1 vssd1 vccd1 vccd1 _13412_/Y sky130_fd_sc_hd__a21oi_1
X_17180_ _17210_/A _17180_/B vssd1 vssd1 vccd1 vccd1 _19411_/D sky130_fd_sc_hd__nor2_1
X_10624_ _18555_/Q _18430_/Q _18039_/Q _18007_/Q _09108_/B _10918_/C1 vssd1 vssd1
+ vccd1 vccd1 _10624_/X sky130_fd_sc_hd__mux4_1
X_14392_ _17699_/A0 _18243_/Q _14412_/S vssd1 vssd1 vccd1 vccd1 _18243_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16131_ _18768_/Q _16141_/B vssd1 vssd1 vccd1 vccd1 _16131_/Y sky130_fd_sc_hd__nand2_1
X_13343_ _17868_/Q _13847_/A2 _13854_/B1 _13342_/X vssd1 vssd1 vccd1 vccd1 _13343_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_194_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10555_ _10850_/A1 _18228_/Q _10634_/S0 _18963_/Q vssd1 vssd1 vccd1 vccd1 _10555_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_183_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16062_ _15845_/A _16069_/A _16059_/X _16061_/X _16048_/A vssd1 vssd1 vccd1 vccd1
+ _18738_/D sky130_fd_sc_hd__a221oi_1
XFILLER_6_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13274_ _15332_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _13274_/Y sky130_fd_sc_hd__nand2_1
XFILLER_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10486_ _10483_/X _10485_/X _10479_/X vssd1 vssd1 vccd1 vccd1 _10486_/Y sky130_fd_sc_hd__a21oi_4
X_15013_ _15013_/A _15013_/B vssd1 vssd1 vccd1 vccd1 _15014_/C sky130_fd_sc_hd__nand2_1
X_12225_ _12241_/A _12225_/B _12226_/B vssd1 vssd1 vccd1 vccd1 _17873_/D sky130_fd_sc_hd__nor3_1
XFILLER_185_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12156_ _17847_/Q _12154_/B _12155_/Y vssd1 vssd1 vccd1 vccd1 _17847_/D sky130_fd_sc_hd__o21a_1
XFILLER_111_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11107_ _11352_/A1 _19635_/Q _18924_/Q _11125_/B2 vssd1 vssd1 vccd1 vccd1 _11107_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16964_ _16964_/A _16964_/B vssd1 vssd1 vccd1 vccd1 _19325_/D sky130_fd_sc_hd__and2_1
X_12087_ _17821_/Q _12087_/B vssd1 vssd1 vccd1 vccd1 _12087_/X sky130_fd_sc_hd__or2_1
XFILLER_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18703_ _18776_/CLK _18703_/D vssd1 vssd1 vccd1 vccd1 _18703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15915_ _18680_/Q _15918_/A2 _15945_/C1 _15914_/X vssd1 vssd1 vccd1 vccd1 _15915_/X
+ sky130_fd_sc_hd__a211o_1
X_11038_ _11428_/A _11037_/X _11508_/B1 vssd1 vssd1 vccd1 vccd1 _11039_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16895_ _19308_/Q _17583_/A _16971_/S vssd1 vssd1 vccd1 vccd1 _16896_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18634_ _19076_/CLK _18634_/D vssd1 vssd1 vccd1 vccd1 _18634_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _18741_/Q _18740_/Q vssd1 vssd1 vccd1 vccd1 _16063_/A sky130_fd_sc_hd__or2_4
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18565_ _19507_/CLK _18565_/D vssd1 vssd1 vccd1 vccd1 _18565_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _13041_/S _12717_/X _12988_/X vssd1 vssd1 vccd1 vccd1 _12989_/Y sky130_fd_sc_hd__o21ai_2
X_15777_ _19486_/Q _19420_/Q vssd1 vssd1 vccd1 vccd1 _15778_/B sky130_fd_sc_hd__or2_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17516_ _18587_/Q _17527_/A1 _17515_/X _17516_/C1 vssd1 vssd1 vccd1 vccd1 _17516_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14728_ input76/X input71/X _14784_/S vssd1 vssd1 vccd1 vccd1 _14728_/X sky130_fd_sc_hd__mux2_8
X_18496_ _18501_/CLK _18496_/D vssd1 vssd1 vccd1 vccd1 _18496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14659_ _16618_/A0 _18465_/Q _14664_/S vssd1 vssd1 vccd1 vccd1 _18465_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17447_ _18112_/Q _17463_/A2 _17445_/X _17446_/X vssd1 vssd1 vccd1 vccd1 _17447_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17378_ _17378_/A _17378_/B vssd1 vssd1 vccd1 vccd1 _19486_/D sky130_fd_sc_hd__and2_1
XFILLER_229_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19117_ _19604_/CLK _19117_/D vssd1 vssd1 vccd1 vccd1 _19117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16329_ _18941_/Q _17661_/A0 _16352_/S vssd1 vssd1 vccd1 vccd1 _18941_/D sky130_fd_sc_hd__mux2_1
XFILLER_229_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19048_ _19075_/CLK _19048_/D vssd1 vssd1 vccd1 vccd1 _19048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput289 _11964_/X vssd1 vssd1 vccd1 vccd1 addr0[4] sky130_fd_sc_hd__buf_4
XFILLER_87_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09703_ _18598_/Q _18169_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09703_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09634_ _09621_/X _09623_/X _10180_/A vssd1 vssd1 vccd1 vccd1 _09634_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_261_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09565_ input111/X input146/X _09651_/S vssd1 vssd1 vccd1 vccd1 _09566_/B sky130_fd_sc_hd__mux2_4
XFILLER_55_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ _11190_/A1 _18139_/Q _18785_/Q _09952_/S _10144_/B1 vssd1 vssd1 vccd1 vccd1
+ _09496_/X sky130_fd_sc_hd__a221o_1
XFILLER_212_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10340_ _10326_/A _10339_/Y _10326_/Y _09611_/A vssd1 vssd1 vccd1 vccd1 _10340_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_279_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10271_ _11488_/A _10271_/B vssd1 vssd1 vccd1 vccd1 _10271_/Y sky130_fd_sc_hd__nor2_1
XFILLER_279_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12010_ _17777_/Q _16611_/A0 _12022_/S vssd1 vssd1 vccd1 vccd1 _17777_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1404 _09539_/S vssd1 vssd1 vccd1 vccd1 _09925_/S sky130_fd_sc_hd__buf_6
XFILLER_155_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1415 _09092_/Y vssd1 vssd1 vccd1 vccd1 fanout1415/X sky130_fd_sc_hd__buf_6
Xfanout1426 _09092_/Y vssd1 vssd1 vccd1 vccd1 _11403_/S sky130_fd_sc_hd__buf_6
XFILLER_24_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1437 _09087_/Y vssd1 vssd1 vccd1 vccd1 _10632_/S sky130_fd_sc_hd__buf_4
XFILLER_94_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1448 _10918_/C1 vssd1 vssd1 vccd1 vccd1 _11559_/S1 sky130_fd_sc_hd__buf_8
XFILLER_266_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1459 _10217_/B vssd1 vssd1 vccd1 vccd1 _10816_/A2 sky130_fd_sc_hd__buf_12
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13961_ _13961_/A _14153_/B vssd1 vssd1 vccd1 vccd1 _13961_/X sky130_fd_sc_hd__or2_1
XFILLER_120_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout494 _14667_/X vssd1 vssd1 vccd1 vccd1 _15001_/A2 sky130_fd_sc_hd__buf_6
XFILLER_86_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15700_ _13818_/A _15111_/A _13838_/X _15112_/B vssd1 vssd1 vccd1 vccd1 _15700_/X
+ sky130_fd_sc_hd__o22a_1
X_12912_ _19427_/Q _12582_/X _12911_/X vssd1 vssd1 vccd1 vccd1 _12912_/X sky130_fd_sc_hd__o21a_2
X_16680_ _19235_/Q _19233_/Q _19232_/Q _16680_/D vssd1 vssd1 vccd1 vccd1 _16690_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_247_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13892_ _13958_/B _14152_/B _13892_/B1 vssd1 vssd1 vccd1 vccd1 _13892_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_73_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15631_ _15631_/A _15631_/B vssd1 vssd1 vccd1 vccd1 _15631_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ _12604_/Y _13312_/A _12842_/X _12841_/X vssd1 vssd1 vccd1 vccd1 _12843_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18350_ _19126_/CLK _18350_/D vssd1 vssd1 vccd1 vccd1 _18350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15562_ _18582_/Q _15581_/C vssd1 vssd1 vccd1 vccd1 _15562_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _19425_/Q _12582_/X _12773_/X vssd1 vssd1 vccd1 vccd1 _12774_/X sky130_fd_sc_hd__o21a_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _19451_/Q _17307_/B vssd1 vssd1 vccd1 vccd1 _17301_/Y sky130_fd_sc_hd__nand2_1
X_14513_ _17715_/A0 _18363_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _18363_/D sky130_fd_sc_hd__mux2_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_48_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19646_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _18777_/Q _11726_/B vssd1 vssd1 vccd1 vccd1 _11725_/X sky130_fd_sc_hd__and2_2
X_18281_ _18741_/CLK _18281_/D vssd1 vssd1 vccd1 vccd1 _18281_/Q sky130_fd_sc_hd__dfxtp_1
X_15493_ _15472_/B _15474_/B _15472_/A vssd1 vssd1 vccd1 vccd1 _15497_/A sky130_fd_sc_hd__a21bo_2
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14444_ _18583_/Q _14452_/B vssd1 vssd1 vccd1 vccd1 _18296_/D sky130_fd_sc_hd__and2_1
X_17232_ _19428_/Q _17241_/B vssd1 vssd1 vccd1 vccd1 _17232_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11656_ _12264_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _12265_/B sky130_fd_sc_hd__and2_4
XFILLER_80_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10607_ _17975_/Q _16820_/A3 _11216_/B1 vssd1 vssd1 vccd1 vccd1 _10607_/X sky130_fd_sc_hd__a21o_1
X_17163_ _17211_/A _17587_/A vssd1 vssd1 vccd1 vccd1 _17462_/A sky130_fd_sc_hd__nand2_1
X_14375_ _18227_/Q _16549_/A0 _14383_/S vssd1 vssd1 vccd1 vccd1 _18227_/D sky130_fd_sc_hd__mux2_1
X_11587_ _11584_/X _11586_/X _11583_/A vssd1 vssd1 vccd1 vccd1 _11587_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16114_ _16078_/X _16113_/Y _12107_/A vssd1 vssd1 vccd1 vccd1 _18759_/D sky130_fd_sc_hd__a21oi_1
XFILLER_183_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13326_ _18113_/Q _13326_/B vssd1 vssd1 vccd1 vccd1 _13327_/B sky130_fd_sc_hd__nor2_1
X_10538_ _19059_/Q _19027_/Q _10613_/S vssd1 vssd1 vccd1 vccd1 _10538_/X sky130_fd_sc_hd__mux2_1
X_17094_ _17181_/B _17116_/A2 _17093_/X _17356_/A vssd1 vssd1 vccd1 vccd1 _19380_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16045_ _18727_/Q _18734_/Q _16051_/S vssd1 vssd1 vccd1 vccd1 _16046_/B sky130_fd_sc_hd__mux2_1
X_13257_ _13257_/A _13257_/B vssd1 vssd1 vccd1 vccd1 _17930_/D sky130_fd_sc_hd__and2_1
X_10469_ _18868_/Q _18900_/Q _10613_/S vssd1 vssd1 vccd1 vccd1 _10469_/X sky130_fd_sc_hd__mux2_1
X_12208_ _17866_/Q _17867_/Q _12208_/C vssd1 vssd1 vccd1 vccd1 _12210_/B sky130_fd_sc_hd__and3_1
XFILLER_124_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13188_ _13188_/A _13188_/B _13188_/C vssd1 vssd1 vccd1 vccd1 _13189_/B sky130_fd_sc_hd__nor3_1
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12139_ _12219_/A _12144_/C vssd1 vssd1 vccd1 vccd1 _12139_/Y sky130_fd_sc_hd__nor2_1
X_17996_ _19630_/CLK _17996_/D vssd1 vssd1 vccd1 vccd1 _17996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16947_ _19321_/Q _17196_/B _16947_/S vssd1 vssd1 vccd1 vccd1 _16948_/B sky130_fd_sc_hd__mux2_1
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16878_ _12492_/A _17928_/Q _16877_/X vssd1 vssd1 vccd1 vccd1 _17575_/A sky130_fd_sc_hd__o21a_4
XFILLER_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18617_ _19641_/CLK _18617_/D vssd1 vssd1 vccd1 vccd1 _18617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15829_ _18621_/Q _17719_/A0 _15829_/S vssd1 vssd1 vccd1 vccd1 _18621_/D sky130_fd_sc_hd__mux2_1
X_19597_ _19629_/CLK _19597_/D vssd1 vssd1 vccd1 vccd1 _19597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09350_ _09348_/X _09349_/X _09350_/S vssd1 vssd1 vccd1 vccd1 _09350_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18548_ _19197_/CLK _18548_/D vssd1 vssd1 vccd1 vccd1 _18548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09281_ _14224_/A _13185_/A vssd1 vssd1 vccd1 vccd1 _09281_/Y sky130_fd_sc_hd__nand2_2
X_18479_ _19320_/CLK _18479_/D vssd1 vssd1 vccd1 vccd1 _18479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08996_ _09028_/B _08996_/B vssd1 vssd1 vccd1 vccd1 _11217_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09617_ _11161_/S _09612_/X _09616_/X vssd1 vssd1 vccd1 vccd1 _09617_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09548_ _09535_/X _09537_/X _10326_/A vssd1 vssd1 vccd1 vccd1 _09548_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09479_ input112/X input147/X _09651_/S vssd1 vssd1 vccd1 vccd1 _09480_/B sky130_fd_sc_hd__mux2_4
XFILLER_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11510_ _18248_/Q _18823_/Q _18451_/Q _18352_/Q _11513_/B2 _11510_/S1 vssd1 vssd1
+ vccd1 vccd1 _11511_/B sky130_fd_sc_hd__mux4_1
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12490_ _12572_/B _12572_/C vssd1 vssd1 vccd1 vccd1 _12553_/C sky130_fd_sc_hd__nand2b_2
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ _18114_/Q _11441_/B vssd1 vssd1 vccd1 vccd1 _11441_/X sky130_fd_sc_hd__or2_2
XFILLER_137_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ _18080_/Q _12461_/A _14340_/A _14159_/Y vssd1 vssd1 vccd1 vccd1 _18080_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11372_ _11219_/A _10163_/B _10757_/B _09039_/B vssd1 vssd1 vccd1 vccd1 _11372_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_192_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ _19335_/Q _13246_/A2 _13246_/B1 _19463_/Q _12570_/C vssd1 vssd1 vccd1 vccd1
+ _13111_/X sky130_fd_sc_hd__a221o_1
XFILLER_124_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10323_ _10323_/A1 _18160_/Q _18806_/Q _10687_/S vssd1 vssd1 vccd1 vccd1 _10323_/X
+ sky130_fd_sc_hd__a22o_1
X_14091_ _17707_/A0 _18031_/Q _14098_/S vssd1 vssd1 vccd1 vccd1 _18031_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_166_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19481_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_152_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13042_ _12895_/Y _13354_/B _13314_/S vssd1 vssd1 vccd1 vccd1 _13042_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10254_ _18161_/Q _11482_/A2 _10253_/X _11406_/B2 vssd1 vssd1 vccd1 vccd1 _10254_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_3_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1201 _12755_/X vssd1 vssd1 vccd1 vccd1 _13912_/A2 sky130_fd_sc_hd__buf_6
X_17850_ _19324_/CLK _17850_/D vssd1 vssd1 vccd1 vccd1 _17850_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1212 _12667_/X vssd1 vssd1 vccd1 vccd1 _14154_/B1 sky130_fd_sc_hd__buf_4
XFILLER_120_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10185_ _10336_/A _10184_/X _11466_/B1 vssd1 vssd1 vccd1 vccd1 _10185_/X sky130_fd_sc_hd__o21a_1
Xfanout1223 _12314_/X vssd1 vssd1 vccd1 vccd1 _13899_/A sky130_fd_sc_hd__buf_4
XFILLER_278_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1234 _12265_/Y vssd1 vssd1 vccd1 vccd1 _12442_/C sky130_fd_sc_hd__buf_6
X_16801_ _19289_/Q _16802_/B vssd1 vssd1 vccd1 vccd1 _16803_/B sky130_fd_sc_hd__nor2_1
Xfanout1245 _08947_/B vssd1 vssd1 vccd1 vccd1 _11451_/B2 sky130_fd_sc_hd__buf_4
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1256 _13807_/A vssd1 vssd1 vccd1 vccd1 _10905_/S sky130_fd_sc_hd__buf_8
X_17781_ _19609_/CLK _17781_/D vssd1 vssd1 vccd1 vccd1 _17781_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1267 _08890_/Y vssd1 vssd1 vccd1 vccd1 _09866_/B sky130_fd_sc_hd__buf_6
Xfanout1278 _11715_/B vssd1 vssd1 vccd1 vccd1 _15006_/B1 sky130_fd_sc_hd__buf_6
X_14993_ _17820_/Q _14992_/X _14993_/S vssd1 vssd1 vccd1 vccd1 _14993_/X sky130_fd_sc_hd__mux2_1
XFILLER_281_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1289 _15037_/S vssd1 vssd1 vccd1 vccd1 _15038_/S sky130_fd_sc_hd__buf_6
XFILLER_47_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19520_ _19552_/CLK _19520_/D vssd1 vssd1 vccd1 vccd1 _19520_/Q sky130_fd_sc_hd__dfxtp_1
X_16732_ _19263_/Q _16734_/C _16731_/X vssd1 vssd1 vccd1 vccd1 _19263_/D sky130_fd_sc_hd__o21ba_1
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13944_ _17854_/Q _13944_/B vssd1 vssd1 vccd1 vccd1 _13944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19451_ _19484_/CLK _19451_/D vssd1 vssd1 vccd1 vccd1 _19451_/Q sky130_fd_sc_hd__dfxtp_1
X_16663_ _19243_/Q _16667_/C vssd1 vssd1 vccd1 vccd1 _16665_/B sky130_fd_sc_hd__nor2_1
X_13875_ _17852_/Q _13942_/A2 _13942_/B1 _17884_/Q vssd1 vssd1 vccd1 vccd1 _13875_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18402_ _19466_/CLK _18402_/D vssd1 vssd1 vccd1 vccd1 _18402_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12826_ _12826_/A vssd1 vssd1 vccd1 vccd1 _12826_/Y sky130_fd_sc_hd__inv_2
X_15614_ _17540_/B1 _15613_/X _15782_/B1 vssd1 vssd1 vccd1 vccd1 _15614_/X sky130_fd_sc_hd__a21o_1
X_19382_ _19483_/CLK _19382_/D vssd1 vssd1 vccd1 vccd1 _19382_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_188_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16594_ _16594_/A0 _19197_/Q _16619_/S vssd1 vssd1 vccd1 vccd1 _19197_/D sky130_fd_sc_hd__mux2_1
X_18333_ _19612_/CLK _18333_/D vssd1 vssd1 vccd1 vccd1 _18333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _19475_/Q _15544_/X _15781_/S vssd1 vssd1 vccd1 vccd1 _15545_/X sky130_fd_sc_hd__mux2_1
X_12757_ _12442_/D _12739_/X _12752_/X _12835_/A vssd1 vssd1 vccd1 vccd1 _12757_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _18516_/Q _18517_/Q _18520_/Q _18519_/Q vssd1 vssd1 vccd1 vccd1 _11708_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_203_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18264_ _19646_/CLK _18264_/D vssd1 vssd1 vccd1 vccd1 _18264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15476_ _15476_/A1 _15475_/X _15499_/B1 vssd1 vssd1 vccd1 vccd1 _15476_/X sky130_fd_sc_hd__a21o_1
X_12688_ _12687_/X _12686_/X _12796_/S vssd1 vssd1 vccd1 vccd1 _12688_/X sky130_fd_sc_hd__mux2_2
XFILLER_129_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14427_ _18566_/Q _14427_/B vssd1 vssd1 vccd1 vccd1 _18279_/D sky130_fd_sc_hd__and2_1
X_17215_ _17556_/A _17120_/Y _17214_/Y _17285_/A vssd1 vssd1 vccd1 vccd1 _17215_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_129_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11639_ _11639_/A _11639_/B vssd1 vssd1 vccd1 vccd1 _13807_/B sky130_fd_sc_hd__xnor2_4
X_18195_ _19628_/CLK _18195_/D vssd1 vssd1 vccd1 vccd1 _18195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14358_ _18210_/Q _16532_/A0 _14377_/S vssd1 vssd1 vccd1 vccd1 _18210_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17146_ _19400_/Q fanout534/X _17433_/A _17212_/B2 vssd1 vssd1 vccd1 vccd1 _17147_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_128_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13309_ _13438_/A _13295_/Y _13563_/B1 vssd1 vssd1 vccd1 vccd1 _13321_/C sky130_fd_sc_hd__a21oi_1
X_17077_ _19372_/Q _17077_/B vssd1 vssd1 vccd1 vccd1 _17077_/X sky130_fd_sc_hd__or2_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14289_ _16607_/A0 _18148_/Q _14301_/S vssd1 vssd1 vccd1 vccd1 _18148_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16028_ _18735_/Q _18727_/Q _16034_/S vssd1 vssd1 vccd1 vccd1 _16028_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08850_ _09494_/A vssd1 vssd1 vccd1 vccd1 _08850_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17979_ _18627_/CLK _17979_/D vssd1 vssd1 vccd1 vccd1 _17979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1790 _10742_/A1 vssd1 vssd1 vccd1 vccd1 _10297_/A1 sky130_fd_sc_hd__buf_6
XFILLER_226_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19649_ _19649_/CLK _19649_/D vssd1 vssd1 vccd1 vccd1 _19649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09402_ _09401_/A _09401_/B _09401_/C vssd1 vssd1 vccd1 vccd1 _09403_/B sky130_fd_sc_hd__o21ai_4
XFILLER_253_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09333_ _17960_/Q _11295_/A2 _08947_/A _17928_/Q _08946_/B vssd1 vssd1 vccd1 vccd1
+ _09333_/Y sky130_fd_sc_hd__a221oi_4
X_09264_ _09262_/X _09263_/X _09264_/S vssd1 vssd1 vccd1 vccd1 _09264_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09195_ _19045_/Q _19013_/Q _10141_/S vssd1 vssd1 vccd1 vccd1 _09195_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08979_ _10419_/S _08979_/B vssd1 vssd1 vccd1 vccd1 _08979_/Y sky130_fd_sc_hd__nand2_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11990_ _14351_/A _14599_/A vssd1 vssd1 vccd1 vccd1 _11990_/Y sky130_fd_sc_hd__nor2_8
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10941_ _11312_/A1 _18152_/Q _18798_/Q _10940_/S vssd1 vssd1 vccd1 vccd1 _10941_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_217_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13660_ _13929_/A1 _13659_/X _13647_/Y vssd1 vssd1 vccd1 vccd1 _13660_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10872_ _11332_/B1 _10870_/X _10871_/X vssd1 vssd1 vccd1 vccd1 _11854_/A sky130_fd_sc_hd__o21ai_1
XFILLER_271_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _13083_/A _13127_/A vssd1 vssd1 vccd1 vccd1 _12615_/A sky130_fd_sc_hd__or2_1
XFILLER_213_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _19380_/Q _13884_/A2 _13589_/X _13590_/X _13884_/C1 vssd1 vssd1 vccd1 vccd1
+ _13591_/X sky130_fd_sc_hd__o221a_4
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15330_/A _15330_/B vssd1 vssd1 vccd1 vccd1 _15330_/Y sky130_fd_sc_hd__nor2_1
X_12542_ _12544_/A _13167_/A vssd1 vssd1 vccd1 vccd1 _12542_/Y sky130_fd_sc_hd__nor2_1
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15261_ _18109_/Q _15132_/X _15260_/X _15382_/B2 vssd1 vssd1 vccd1 vccd1 _15262_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_12473_ _12507_/A _12514_/A vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__nand2_8
XFILLER_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17000_ _17575_/A _17008_/A2 _16999_/X _17559_/A vssd1 vssd1 vccd1 vccd1 _19336_/D
+ sky130_fd_sc_hd__o211a_1
X_14212_ _18104_/Q _14244_/B vssd1 vssd1 vccd1 vccd1 _14212_/X sky130_fd_sc_hd__or2_1
X_11424_ _09967_/S _11419_/X _11423_/X vssd1 vssd1 vccd1 vccd1 _11424_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15192_ _17219_/A _15192_/B _15192_/C vssd1 vssd1 vccd1 vccd1 _15192_/Y sky130_fd_sc_hd__nor3_1
XANTENNA_8 _18275_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _14143_/A _14143_/B _14143_/C _13149_/X vssd1 vssd1 vccd1 vccd1 _14144_/A
+ sky130_fd_sc_hd__or4b_2
X_11355_ _11355_/A1 _11354_/X _11623_/A1 vssd1 vssd1 vccd1 vccd1 _11356_/B sky130_fd_sc_hd__a21o_1
XFILLER_193_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _10307_/A _12658_/B vssd1 vssd1 vccd1 vccd1 _11636_/A sky130_fd_sc_hd__or2_4
X_18951_ _19612_/CLK _18951_/D vssd1 vssd1 vccd1 vccd1 _18951_/Q sky130_fd_sc_hd__dfxtp_1
X_14074_ _16459_/B _14074_/B _14074_/C vssd1 vssd1 vccd1 vccd1 _16426_/A sky130_fd_sc_hd__and3b_4
XFILLER_4_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11286_ _10745_/S _11285_/X _11286_/B1 vssd1 vssd1 vccd1 vccd1 _11286_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_112_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17902_ _18201_/CLK _17902_/D vssd1 vssd1 vccd1 vccd1 _17902_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_140_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13025_ _13929_/A1 _13024_/X _13008_/Y vssd1 vssd1 vccd1 vccd1 _13027_/B sky130_fd_sc_hd__a21o_1
XFILLER_279_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10237_ _11064_/B1 _10235_/Y _10236_/X vssd1 vssd1 vccd1 vccd1 _10237_/X sky130_fd_sc_hd__o21a_1
X_18882_ _19614_/CLK _18882_/D vssd1 vssd1 vccd1 vccd1 _18882_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1020 _14973_/A1 vssd1 vssd1 vccd1 vccd1 _14912_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_266_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1031 _16597_/A0 vssd1 vssd1 vccd1 vccd1 _17697_/A0 sky130_fd_sc_hd__clkbuf_4
X_17833_ _17865_/CLK _17833_/D vssd1 vssd1 vccd1 vccd1 _17833_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1042 _09140_/S vssd1 vssd1 vccd1 vccd1 _09643_/A sky130_fd_sc_hd__buf_4
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10168_ _18468_/Q _18369_/Q _10168_/S vssd1 vssd1 vccd1 vccd1 _10168_/X sky130_fd_sc_hd__mux2_1
Xfanout1053 _17603_/B1 vssd1 vssd1 vccd1 vccd1 _17588_/B1 sky130_fd_sc_hd__buf_6
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1064 _13486_/A1 vssd1 vssd1 vccd1 vccd1 _13958_/B sky130_fd_sc_hd__buf_6
XFILLER_282_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1075 _12460_/Y vssd1 vssd1 vccd1 vccd1 _14027_/A2 sky130_fd_sc_hd__buf_4
XFILLER_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1086 _16462_/A0 vssd1 vssd1 vccd1 vccd1 _17661_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_281_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17764_ _19201_/CLK _17764_/D vssd1 vssd1 vccd1 vccd1 _17764_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1097 _09055_/X vssd1 vssd1 vccd1 vccd1 _11624_/A1 sky130_fd_sc_hd__buf_8
X_10099_ _18624_/Q _18195_/Q _10099_/S vssd1 vssd1 vccd1 vccd1 _10099_/X sky130_fd_sc_hd__mux2_1
X_14976_ _14996_/A1 _14975_/X _15006_/B1 vssd1 vssd1 vccd1 vccd1 _14976_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_208_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19503_ _19552_/CLK _19503_/D vssd1 vssd1 vccd1 vccd1 _19503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19213_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16715_ _19258_/Q _16715_/B vssd1 vssd1 vccd1 vccd1 _16722_/C sky130_fd_sc_hd__and2_1
X_13927_ _17853_/Q _13944_/B _13920_/X _13926_/X vssd1 vssd1 vccd1 vccd1 _13927_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_228_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17695_ _17695_/A0 _19621_/Q _17718_/S vssd1 vssd1 vccd1 vccd1 _19621_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19434_ _19530_/CLK _19434_/D vssd1 vssd1 vccd1 vccd1 _19434_/Q sky130_fd_sc_hd__dfxtp_1
X_16646_ _19238_/Q _16649_/C vssd1 vssd1 vccd1 vccd1 _16648_/A sky130_fd_sc_hd__and2_1
XFILLER_228_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _13758_/A _13843_/Y _13956_/B1 vssd1 vssd1 vccd1 vccd1 _13858_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_211_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19365_ _19458_/CLK _19365_/D vssd1 vssd1 vccd1 vccd1 _19365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12809_ _12708_/X _12704_/X _12813_/S vssd1 vssd1 vccd1 vccd1 _12810_/A sky130_fd_sc_hd__mux2_1
X_16577_ _16610_/A0 _19181_/Q _16589_/S vssd1 vssd1 vccd1 vccd1 _19181_/D sky130_fd_sc_hd__mux2_1
XFILLER_210_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13789_ _13637_/A _14026_/B _13775_/X vssd1 vssd1 vccd1 vccd1 _13791_/B sky130_fd_sc_hd__o21ai_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18316_ _19595_/CLK _18316_/D vssd1 vssd1 vccd1 vccd1 _18316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ _18120_/Q _15133_/Y _15527_/X _15452_/A vssd1 vssd1 vccd1 vccd1 _15531_/A
+ sky130_fd_sc_hd__a22o_1
X_19296_ _19304_/CLK _19296_/D vssd1 vssd1 vccd1 vccd1 _19296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18247_ _18884_/CLK _18247_/D vssd1 vssd1 vccd1 vccd1 _18247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15459_ _15385_/A _15386_/Y _15456_/C _15456_/D _15384_/Y vssd1 vssd1 vccd1 vccd1
+ _15459_/X sky130_fd_sc_hd__a2111o_2
XFILLER_128_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18178_ _19630_/CLK _18178_/D vssd1 vssd1 vccd1 vccd1 _18178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17129_ _17129_/A _17565_/B vssd1 vssd1 vccd1 vccd1 _17129_/Y sky130_fd_sc_hd__nor2_2
XFILLER_274_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09951_ _18237_/Q _18812_/Q _09952_/S vssd1 vssd1 vccd1 vccd1 _09951_/X sky130_fd_sc_hd__mux2_1
X_08902_ _09494_/A _12024_/A vssd1 vssd1 vccd1 vccd1 _08902_/Y sky130_fd_sc_hd__nand2_2
XFILLER_258_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _18018_/Q _17986_/Q _10054_/S vssd1 vssd1 vccd1 vccd1 _09882_/X sky130_fd_sc_hd__mux2_1
XFILLER_253_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08833_ _18110_/Q vssd1 vssd1 vccd1 vccd1 _14224_/A sky130_fd_sc_hd__inv_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_409 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09316_ _12600_/A _09317_/B vssd1 vssd1 vccd1 vccd1 _13195_/S sky130_fd_sc_hd__or2_2
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09247_ _17961_/Q _11295_/A2 _08947_/A _17929_/Q _08946_/B vssd1 vssd1 vccd1 vccd1
+ _09247_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_194_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09178_ _09176_/X _09177_/X _10169_/S vssd1 vssd1 vccd1 vccd1 _09178_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11140_ _13485_/A vssd1 vssd1 vccd1 vccd1 _11676_/A sky130_fd_sc_hd__inv_2
XFILLER_134_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11071_ _11562_/S _11070_/X _11069_/X _11084_/S vssd1 vssd1 vccd1 vccd1 _11071_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput101 dout0[62] vssd1 vssd1 vccd1 vccd1 input101/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput112 dout1[14] vssd1 vssd1 vccd1 vccd1 input112/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10022_ _11252_/S _10021_/X _10016_/X _09107_/D vssd1 vssd1 vccd1 vccd1 _10022_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput123 dout1[24] vssd1 vssd1 vccd1 vccd1 input123/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput134 dout1[34] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__buf_2
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 dout1[44] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_hd__clkbuf_2
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput156 dout1[54] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__buf_2
XFILLER_237_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput167 dout1[6] vssd1 vssd1 vccd1 vccd1 input167/X sky130_fd_sc_hd__clkbuf_2
X_14830_ _12053_/A _14829_/X _14993_/S vssd1 vssd1 vccd1 vccd1 _14830_/X sky130_fd_sc_hd__mux2_1
XFILLER_263_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput178 irq[1] vssd1 vssd1 vccd1 vccd1 input178/X sky130_fd_sc_hd__clkbuf_4
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 jtag_tms vssd1 vssd1 vccd1 vccd1 _16075_/A sky130_fd_sc_hd__buf_6
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ _14759_/X _14760_/X _14913_/B1 vssd1 vssd1 vccd1 vccd1 _14761_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11973_ _18737_/Q _18734_/Q _18733_/Q _18735_/Q vssd1 vssd1 vccd1 vccd1 _11973_/X
+ sky130_fd_sc_hd__or4b_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16500_ _16500_/A0 _19106_/Q _16521_/S vssd1 vssd1 vccd1 vccd1 _19106_/D sky130_fd_sc_hd__mux2_1
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _17847_/Q _13744_/A2 _13744_/B1 _17879_/Q vssd1 vssd1 vccd1 vccd1 _13712_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ _11311_/C1 _10923_/X _10922_/X _10930_/S vssd1 vssd1 vccd1 vccd1 _10924_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_260_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _12276_/B _14692_/A2 _15834_/C vssd1 vssd1 vccd1 vccd1 _14692_/X sky130_fd_sc_hd__o21ba_1
X_17480_ _13545_/B _17520_/A2 _17532_/A2 _17808_/Q _17538_/A vssd1 vssd1 vccd1 vccd1
+ _17480_/X sky130_fd_sc_hd__a221o_1
XFILLER_232_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ _19039_/Q _16431_/A1 _16454_/S vssd1 vssd1 vccd1 vccd1 _19039_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13643_ _13704_/C _13643_/B vssd1 vssd1 vccd1 vccd1 _13643_/X sky130_fd_sc_hd__or2_2
X_10855_ _19055_/Q _19023_/Q _10864_/S vssd1 vssd1 vccd1 vccd1 _10855_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19150_ _19226_/CLK _19150_/D vssd1 vssd1 vccd1 vccd1 _19150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13574_ _13968_/B2 _13573_/X _13565_/Y vssd1 vssd1 vccd1 vccd1 _13574_/X sky130_fd_sc_hd__a21o_1
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _16462_/A0 _18973_/Q _16385_/S vssd1 vssd1 vccd1 vccd1 _18973_/D sky130_fd_sc_hd__mux2_1
X_10786_ _18647_/Q _18069_/Q _19088_/Q _18992_/Q _11302_/S _11559_/S1 vssd1 vssd1
+ vccd1 vccd1 _10786_/X sky130_fd_sc_hd__mux4_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18101_ _18593_/CLK _18101_/D vssd1 vssd1 vccd1 vccd1 _18101_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12525_ _13167_/A _12768_/B _12577_/B vssd1 vssd1 vccd1 vccd1 _12525_/X sky130_fd_sc_hd__a21o_1
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15313_ _15313_/A _15313_/B vssd1 vssd1 vccd1 vccd1 _15313_/Y sky130_fd_sc_hd__nand2_1
XFILLER_184_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16293_ _17625_/A _17691_/B vssd1 vssd1 vccd1 vccd1 _16293_/Y sky130_fd_sc_hd__nand2_2
X_19081_ _19118_/CLK _19081_/D vssd1 vssd1 vccd1 vccd1 _19081_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_181_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18279_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18032_ _19586_/CLK _18032_/D vssd1 vssd1 vccd1 vccd1 _18032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12456_ _16819_/A _16819_/B _16836_/S vssd1 vssd1 vccd1 vccd1 _14669_/B sky130_fd_sc_hd__o21ai_2
X_15244_ _15220_/Y _15222_/B _15218_/Y vssd1 vssd1 vccd1 vccd1 _15248_/B sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_110_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19273_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11407_ _11380_/X _11383_/X _11484_/B1 vssd1 vssd1 vccd1 vccd1 _11407_/X sky130_fd_sc_hd__a21o_1
X_15175_ _14214_/A _15132_/X _15174_/Y _12318_/A vssd1 vssd1 vccd1 vccd1 _15177_/B
+ sky130_fd_sc_hd__o22a_1
X_12387_ _12420_/A1 _12409_/A2 _09323_/X _12417_/B1 _18389_/Q vssd1 vssd1 vccd1 vccd1
+ _12388_/B sky130_fd_sc_hd__o32ai_2
XFILLER_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14126_ _16543_/A0 _18065_/Q _14140_/S vssd1 vssd1 vccd1 vccd1 _18065_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ _18546_/Q _18421_/Q _18030_/Q _17998_/Q _11353_/B2 _11338_/S1 vssd1 vssd1
+ vccd1 vccd1 _11338_/X sky130_fd_sc_hd__mux4_1
XFILLER_259_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18934_ _19645_/CLK _18934_/D vssd1 vssd1 vccd1 vccd1 _18934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14057_ _16607_/A0 _17999_/Q _14064_/S vssd1 vssd1 vccd1 vccd1 _17999_/D sky130_fd_sc_hd__mux2_1
X_11269_ _11277_/A1 _18148_/Q _18794_/Q _10744_/S vssd1 vssd1 vccd1 vccd1 _11269_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13008_ _15194_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _13008_/Y sky130_fd_sc_hd__nor2_1
X_18865_ _19601_/CLK _18865_/D vssd1 vssd1 vccd1 vccd1 _18865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17816_ _19492_/CLK _17816_/D vssd1 vssd1 vccd1 vccd1 _17816_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_283_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18796_ _19635_/CLK _18796_/D vssd1 vssd1 vccd1 vccd1 _18796_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17747_ _18647_/Q vssd1 vssd1 vccd1 vccd1 _18647_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_282_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14959_ _14979_/A1 _18272_/Q _14958_/Y _11712_/A vssd1 vssd1 vccd1 vccd1 _14959_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17678_ _17678_/A0 _19605_/Q _17690_/S vssd1 vssd1 vccd1 vccd1 _19605_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19417_ _19482_/CLK _19417_/D vssd1 vssd1 vccd1 vccd1 _19417_/Q sky130_fd_sc_hd__dfxtp_1
X_16629_ _12312_/B _16628_/X _17725_/C1 vssd1 vssd1 vccd1 vccd1 _19231_/D sky130_fd_sc_hd__a21oi_1
XFILLER_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19348_ _19485_/CLK _19348_/D vssd1 vssd1 vccd1 vccd1 _19348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09101_ _14350_/A _09857_/A1 _09099_/Y _16392_/C _09097_/Y vssd1 vssd1 vccd1 vccd1
+ _09101_/X sky130_fd_sc_hd__o221a_1
XFILLER_241_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19279_ _19280_/CLK _19279_/D vssd1 vssd1 vccd1 vccd1 _19279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09032_ _09043_/A _09032_/B vssd1 vssd1 vccd1 vccd1 _09325_/C sky130_fd_sc_hd__nand2_1
XFILLER_163_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout802 _16189_/S vssd1 vssd1 vccd1 vccd1 _16192_/S sky130_fd_sc_hd__buf_12
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09934_ _09932_/X _09933_/X _10265_/A vssd1 vssd1 vccd1 vccd1 _09935_/B sky130_fd_sc_hd__mux2_1
Xfanout813 _14377_/S vssd1 vssd1 vccd1 vccd1 _14383_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_277_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout824 _14273_/Y vssd1 vssd1 vccd1 vccd1 _14277_/S sky130_fd_sc_hd__buf_12
Xfanout835 _16543_/A0 vssd1 vssd1 vccd1 vccd1 _17676_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout846 _16314_/A0 vssd1 vssd1 vccd1 vccd1 _17712_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout857 _10713_/A2 vssd1 vssd1 vccd1 vccd1 _16548_/A0 sky130_fd_sc_hd__clkbuf_4
X_09865_ _09862_/X _09863_/Y _09141_/A vssd1 vssd1 vccd1 vccd1 _09898_/A sky130_fd_sc_hd__a21o_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout868 _10312_/X vssd1 vssd1 vccd1 vccd1 _10341_/A2 sky130_fd_sc_hd__clkbuf_16
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout879 _15832_/A1 vssd1 vssd1 vccd1 vccd1 _16490_/A0 sky130_fd_sc_hd__clkbuf_4
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08816_ _08816_/A vssd1 vssd1 vccd1 vccd1 _12089_/A sky130_fd_sc_hd__inv_6
XFILLER_100_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _08874_/D _09795_/X _11286_/B1 vssd1 vssd1 vccd1 vccd1 _09796_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_206 _18572_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_217 _17913_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 _18386_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_239 _18395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _09777_/A _11490_/B _10639_/X vssd1 vssd1 vccd1 vccd1 _10677_/A sky130_fd_sc_hd__o21ai_4
XFILLER_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10571_ _18650_/Q _10645_/S vssd1 vssd1 vccd1 vccd1 _10571_/X sky130_fd_sc_hd__or2_1
XFILLER_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12310_ _14671_/A _12308_/X _16836_/S vssd1 vssd1 vccd1 vccd1 _12311_/A sky130_fd_sc_hd__o21ai_2
XFILLER_182_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13290_ _13936_/B2 _13273_/Y _13287_/Y _13289_/Y _13185_/A vssd1 vssd1 vccd1 vccd1
+ _13290_/X sky130_fd_sc_hd__a221o_1
XFILLER_213_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12241_ _12241_/A _12241_/B _12242_/B vssd1 vssd1 vccd1 vccd1 _17879_/D sky130_fd_sc_hd__nor3_1
XFILLER_6_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12172_ _17853_/Q _12170_/B _12171_/Y vssd1 vssd1 vccd1 vccd1 _17853_/D sky130_fd_sc_hd__o21a_1
XFILLER_162_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11123_ _10040_/S _11120_/X _11122_/X vssd1 vssd1 vccd1 vccd1 _11131_/B sky130_fd_sc_hd__a21oi_1
X_16980_ _17555_/B _17217_/B vssd1 vssd1 vccd1 vccd1 _16980_/X sky130_fd_sc_hd__or2_4
XFILLER_3_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15931_ _18686_/Q _15943_/A2 _15930_/X _16764_/B1 vssd1 vssd1 vccd1 vccd1 _18686_/D
+ sky130_fd_sc_hd__o211a_1
X_11054_ _11039_/Y _11052_/X _11053_/X vssd1 vssd1 vccd1 vccd1 _11054_/X sky130_fd_sc_hd__o21a_4
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10005_ _17984_/Q _11224_/B _09996_/X _11569_/S1 vssd1 vssd1 vccd1 vccd1 _10005_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _19620_/CLK _18650_/D vssd1 vssd1 vccd1 vccd1 _18650_/Q sky130_fd_sc_hd__dfxtp_4
X_15862_ _18663_/Q _15949_/A2 _15860_/X _15861_/X _15910_/C1 vssd1 vssd1 vccd1 vccd1
+ _18663_/D sky130_fd_sc_hd__o221a_1
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17601_ _15093_/A _17592_/X _17623_/B1 vssd1 vssd1 vccd1 vccd1 _17601_/X sky130_fd_sc_hd__a21o_1
XFILLER_76_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ _15006_/A1 _14812_/X _14875_/B1 vssd1 vssd1 vccd1 vccd1 _14813_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _19444_/CLK _18581_/D vssd1 vssd1 vccd1 vccd1 _18581_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_264_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _19455_/Q _15793_/A2 _17208_/A vssd1 vssd1 vccd1 vccd1 _15793_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17532_ _17818_/Q _17532_/A2 _17538_/A _17531_/Y vssd1 vssd1 vccd1 vccd1 _17532_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _18106_/Q _14801_/B _14690_/Y _14743_/X vssd1 vssd1 vccd1 vccd1 _14744_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_217_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11956_ _11666_/A _11777_/Y _11663_/A vssd1 vssd1 vccd1 vccd1 _14344_/C sky130_fd_sc_hd__a21o_1
XFILLER_233_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ _12641_/A _10908_/B vssd1 vssd1 vccd1 vccd1 _13600_/S sky130_fd_sc_hd__and2_4
XFILLER_83_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17463_ _18115_/Q _17463_/A2 _17461_/X _17462_/Y vssd1 vssd1 vccd1 vccd1 _17463_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_205_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14675_ _14675_/A _14675_/B _14675_/C vssd1 vssd1 vccd1 vccd1 _14688_/C sky130_fd_sc_hd__or3_4
X_11887_ _10342_/B _11845_/B _11887_/B1 vssd1 vssd1 vccd1 vccd1 _11890_/B sky130_fd_sc_hd__o21ai_2
XFILLER_233_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19202_ _19625_/CLK _19202_/D vssd1 vssd1 vccd1 vccd1 _19202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16414_ _17712_/A0 _19023_/Q _16420_/S vssd1 vssd1 vccd1 vccd1 _19023_/D sky130_fd_sc_hd__mux2_1
X_13626_ _17844_/Q _13846_/B vssd1 vssd1 vccd1 vccd1 _13626_/Y sky130_fd_sc_hd__nor2_1
X_10838_ _18991_/Q _10838_/B vssd1 vssd1 vccd1 vccd1 _10838_/X sky130_fd_sc_hd__or2_1
X_17394_ _17394_/A _17423_/B vssd1 vssd1 vccd1 vccd1 _17394_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ _19133_/CLK _19133_/D vssd1 vssd1 vccd1 vccd1 _19133_/Q sky130_fd_sc_hd__dfxtp_1
X_16345_ _18957_/Q _17644_/A0 _16355_/S vssd1 vssd1 vccd1 vccd1 _18957_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10769_ _18615_/Q _18186_/Q _11576_/S vssd1 vssd1 vccd1 vccd1 _10769_/X sky130_fd_sc_hd__mux2_1
X_13557_ _19347_/Q _13883_/A2 _13883_/B1 _19475_/Q _13883_/C1 vssd1 vssd1 vccd1 vccd1
+ _13557_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19064_ _19647_/CLK _19064_/D vssd1 vssd1 vccd1 vccd1 _19064_/Q sky130_fd_sc_hd__dfxtp_1
X_12508_ _12851_/B _12576_/A vssd1 vssd1 vccd1 vccd1 _12579_/A sky130_fd_sc_hd__or2_4
XFILLER_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13488_ _13962_/B _13487_/X _11139_/B vssd1 vssd1 vccd1 vccd1 _13488_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16276_ _17641_/A0 _18890_/Q _16278_/S vssd1 vssd1 vccd1 vccd1 _18890_/D sky130_fd_sc_hd__mux2_1
XFILLER_218_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18015_ _19134_/CLK _18015_/D vssd1 vssd1 vccd1 vccd1 _18015_/Q sky130_fd_sc_hd__dfxtp_1
X_12439_ _12439_/A _12443_/C vssd1 vssd1 vccd1 vccd1 _12762_/A sky130_fd_sc_hd__nor2_4
X_15227_ _19430_/Q _15411_/B _15731_/B1 _15226_/X vssd1 vssd1 vccd1 vccd1 _15236_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_218_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput405 _11927_/X vssd1 vssd1 vccd1 vccd1 din0[7] sky130_fd_sc_hd__buf_4
Xoutput416 _18486_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[15] sky130_fd_sc_hd__buf_4
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput427 _18496_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[25] sky130_fd_sc_hd__buf_4
Xoutput438 _18477_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[6] sky130_fd_sc_hd__buf_4
XFILLER_154_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15158_ _15137_/A _15137_/B _15157_/X vssd1 vssd1 vccd1 vccd1 _15171_/B sky130_fd_sc_hd__a21o_1
Xoutput449 _18737_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[4] sky130_fd_sc_hd__buf_4
XFILLER_99_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14109_ _16526_/A0 _18048_/Q _14131_/S vssd1 vssd1 vccd1 vccd1 _18048_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15089_ _19388_/Q _15092_/B _15089_/C vssd1 vssd1 vccd1 vccd1 _15093_/B sky130_fd_sc_hd__and3_1
XFILLER_102_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18917_ _19628_/CLK _18917_/D vssd1 vssd1 vccd1 vccd1 _18917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09650_ _09012_/A _09907_/A _09649_/X _09650_/B1 _18377_/Q vssd1 vssd1 vccd1 vccd1
+ _09650_/X sky130_fd_sc_hd__o32a_1
XFILLER_227_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18848_ _18880_/CLK _18848_/D vssd1 vssd1 vccd1 vccd1 _18848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09581_ _18599_/Q _18170_/Q _10362_/S vssd1 vssd1 vccd1 vccd1 _09581_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18779_ _18875_/CLK _18779_/D vssd1 vssd1 vccd1 vccd1 _18779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_283_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09015_ _18380_/Q _09650_/B1 _10085_/A vssd1 vssd1 vccd1 vccd1 _09015_/X sky130_fd_sc_hd__o21a_1
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1608 _15103_/Y vssd1 vssd1 vccd1 vccd1 _17527_/A1 sky130_fd_sc_hd__buf_4
Xfanout610 _11887_/B1 vssd1 vssd1 vccd1 vccd1 _11952_/A2 sky130_fd_sc_hd__buf_12
XFILLER_120_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout621 _17118_/X vssd1 vssd1 vccd1 vccd1 _17158_/B2 sky130_fd_sc_hd__buf_6
Xfanout1619 _09010_/Y vssd1 vssd1 vccd1 vccd1 _09991_/A sky130_fd_sc_hd__buf_6
XFILLER_259_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09917_ _18627_/Q _18049_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _09917_/X sky130_fd_sc_hd__mux2_1
Xfanout632 _12744_/Y vssd1 vssd1 vccd1 vccd1 _13413_/B1 sky130_fd_sc_hd__buf_2
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout643 _17050_/X vssd1 vssd1 vccd1 vccd1 _17108_/A2 sky130_fd_sc_hd__buf_6
Xfanout654 _13921_/S vssd1 vssd1 vccd1 vccd1 _13946_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout665 _12570_/A vssd1 vssd1 vccd1 vccd1 _13654_/A2 sky130_fd_sc_hd__buf_4
XFILLER_101_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout676 _13950_/B1 vssd1 vssd1 vccd1 vccd1 _13883_/B1 sky130_fd_sc_hd__buf_6
XFILLER_274_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout687 _12559_/X vssd1 vssd1 vccd1 vccd1 _12560_/B sky130_fd_sc_hd__buf_6
XFILLER_101_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09848_ _10707_/A _09843_/X _09847_/X _09534_/S vssd1 vssd1 vccd1 vccd1 _09848_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_258_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout698 _12545_/Y vssd1 vssd1 vccd1 vccd1 _13625_/B1 sky130_fd_sc_hd__buf_2
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09776_/X _09777_/Y _09946_/B1 vssd1 vssd1 vccd1 vccd1 _09779_/X sky130_fd_sc_hd__a21o_1
XFILLER_234_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11810_/A _11818_/B _11810_/C vssd1 vssd1 vccd1 vccd1 _11810_/X sky130_fd_sc_hd__and3_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12790_/A vssd1 vssd1 vccd1 vccd1 _12790_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _18567_/Q _11741_/A2 _11799_/B _11740_/Y vssd1 vssd1 vccd1 vccd1 _11741_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14460_ _18312_/Q _17664_/A0 _14483_/S vssd1 vssd1 vccd1 vccd1 _18312_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11672_ _13597_/A _11672_/B vssd1 vssd1 vccd1 vccd1 _13611_/B sky130_fd_sc_hd__xnor2_4
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10623_ _10623_/A _10623_/B vssd1 vssd1 vccd1 vccd1 _10623_/Y sky130_fd_sc_hd__nand2_1
X_13411_ _13411_/A _13411_/B vssd1 vssd1 vccd1 vccd1 _14147_/A sky130_fd_sc_hd__xnor2_2
XFILLER_186_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14391_ _17698_/A0 _18242_/Q _14412_/S vssd1 vssd1 vccd1 vccd1 _18242_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16130_ _16140_/A1 _16129_/Y _16142_/B1 vssd1 vssd1 vccd1 vccd1 _18767_/D sky130_fd_sc_hd__a21oi_1
X_13342_ _19309_/Q _12583_/Y _13340_/X _13341_/X vssd1 vssd1 vccd1 vccd1 _13342_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_195_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ _10618_/S _10549_/X _10553_/X vssd1 vssd1 vccd1 vccd1 _10554_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_183_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16061_ _16034_/S _16063_/B _16075_/B _16020_/A vssd1 vssd1 vccd1 vccd1 _16061_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13273_ _13326_/B _13273_/B vssd1 vssd1 vccd1 vccd1 _13273_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10485_ _10841_/C1 _10484_/X _09106_/B vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12224_ _17872_/Q _17873_/Q _12224_/C vssd1 vssd1 vccd1 vccd1 _12226_/B sky130_fd_sc_hd__and3_1
X_15012_ _08830_/Y _14666_/X _12271_/A _17159_/A vssd1 vssd1 vccd1 vccd1 _18503_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_182_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12155_ _12241_/A _12160_/C vssd1 vssd1 vccd1 vccd1 _12155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11106_ _11611_/S _11106_/B vssd1 vssd1 vccd1 vccd1 _11106_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16963_ _19325_/Q _17208_/B _16963_/S vssd1 vssd1 vccd1 vccd1 _16964_/B sky130_fd_sc_hd__mux2_1
X_12086_ _12442_/A _12086_/A2 _12085_/X _17419_/C1 vssd1 vssd1 vccd1 vccd1 _17820_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18702_ _18776_/CLK _18702_/D vssd1 vssd1 vccd1 vccd1 _18702_/Q sky130_fd_sc_hd__dfxtp_1
X_15914_ _15914_/A _15947_/S _15923_/C vssd1 vssd1 vccd1 vccd1 _15914_/X sky130_fd_sc_hd__and3_1
X_11037_ _11035_/X _11036_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _11037_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16894_ _16970_/A1 _17932_/Q _16893_/X vssd1 vssd1 vccd1 vccd1 _17583_/A sky130_fd_sc_hd__o21a_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18633_ _19591_/CLK _18633_/D vssd1 vssd1 vccd1 vccd1 _18633_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_280_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _15845_/A _15845_/B vssd1 vssd1 vccd1 vccd1 _15853_/A sky130_fd_sc_hd__nor2_8
XFILLER_92_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18564_ _19492_/CLK _18564_/D vssd1 vssd1 vccd1 vccd1 _18564_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _19486_/Q _19420_/Q vssd1 vssd1 vccd1 vccd1 _15776_/X sky130_fd_sc_hd__and2_1
XFILLER_92_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _13089_/A _12988_/B vssd1 vssd1 vccd1 vccd1 _12988_/X sky130_fd_sc_hd__or2_2
XFILLER_220_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _11641_/Y _17520_/A2 _17532_/A2 _17815_/Q _17538_/A vssd1 vssd1 vccd1 vccd1
+ _17515_/X sky130_fd_sc_hd__a221o_1
X_14727_ _14865_/A1 _14725_/X _14875_/B1 vssd1 vssd1 vccd1 vccd1 _14727_/Y sky130_fd_sc_hd__o21ai_2
X_18495_ _18501_/CLK _18495_/D vssd1 vssd1 vccd1 vccd1 _18495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11939_ _11939_/A1 _11853_/B _11945_/B1 input225/X vssd1 vssd1 vccd1 vccd1 _11939_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_233_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17446_ _18573_/Q _15103_/Y _17546_/A2 vssd1 vssd1 vccd1 vccd1 _17446_/X sky130_fd_sc_hd__o21a_1
XFILLER_221_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14658_ _17717_/A0 _18464_/Q _14664_/S vssd1 vssd1 vccd1 vccd1 _18464_/D sky130_fd_sc_hd__mux2_1
XFILLER_221_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13609_ _15481_/B _13605_/X _13608_/X _13869_/B2 vssd1 vssd1 vccd1 vccd1 _13610_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_220_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17377_ _19486_/Q _17211_/B _17377_/S vssd1 vssd1 vccd1 vccd1 _17378_/B sky130_fd_sc_hd__mux2_1
X_14589_ _18403_/Q _14589_/A2 _14589_/B1 input33/X vssd1 vssd1 vccd1 vccd1 _14590_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_174_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19116_ _19148_/CLK _19116_/D vssd1 vssd1 vccd1 vccd1 _19116_/Q sky130_fd_sc_hd__dfxtp_1
X_16328_ _18940_/Q _16461_/A0 _16355_/S vssd1 vssd1 vccd1 vccd1 _18940_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19047_ _19047_/CLK _19047_/D vssd1 vssd1 vccd1 vccd1 _19047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16259_ _16292_/A0 _18874_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _18874_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09702_ _18240_/Q _18815_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__mux2_1
XFILLER_261_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09633_ _11173_/S _09632_/X _09631_/X vssd1 vssd1 vccd1 vccd1 _09633_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09564_ _11691_/B1 _09991_/A _09563_/X _11692_/A1 _18378_/Q vssd1 vssd1 vccd1 vccd1
+ _09564_/X sky130_fd_sc_hd__o32a_1
XFILLER_64_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09495_ _18849_/Q _10364_/B _09494_/X _12389_/A1 vssd1 vssd1 vccd1 vccd1 _09495_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_169_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10270_ _10239_/A _10269_/X _10239_/Y _11790_/B vssd1 vssd1 vccd1 vccd1 _10271_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_105_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1405 _09539_/S vssd1 vssd1 vccd1 vccd1 _11472_/C sky130_fd_sc_hd__buf_2
XFILLER_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1416 _11481_/C vssd1 vssd1 vccd1 vccd1 _11395_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_78_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1427 _09137_/S vssd1 vssd1 vccd1 vccd1 _09107_/D sky130_fd_sc_hd__buf_12
XFILLER_132_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1438 _09534_/S vssd1 vssd1 vccd1 vccd1 _11567_/S sky130_fd_sc_hd__buf_6
XFILLER_259_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1449 _09086_/Y vssd1 vssd1 vccd1 vccd1 _10918_/C1 sky130_fd_sc_hd__buf_6
XFILLER_150_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13960_ _11627_/Y _12663_/B _13959_/X vssd1 vssd1 vccd1 vccd1 _14153_/B sky130_fd_sc_hd__o21ai_4
XFILLER_280_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout495 _11949_/B1 vssd1 vssd1 vccd1 vccd1 _11935_/B1 sky130_fd_sc_hd__buf_6
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12911_ _19395_/Q _12579_/Y _12771_/X _12910_/X _12581_/Y vssd1 vssd1 vccd1 vccd1
+ _12911_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13891_ _13891_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _14152_/B sky130_fd_sc_hd__xnor2_4
XFILLER_111_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15630_ _15628_/X _15630_/B vssd1 vssd1 vccd1 vccd1 _15631_/B sky130_fd_sc_hd__nand2b_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _12842_/A _12842_/B vssd1 vssd1 vccd1 vccd1 _12842_/X sky130_fd_sc_hd__or2_1
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _18582_/Q _18581_/Q _15561_/C vssd1 vssd1 vccd1 vccd1 _15561_/X sky130_fd_sc_hd__and3_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _19393_/Q _12579_/Y _12771_/X _12772_/X _12581_/Y vssd1 vssd1 vccd1 vccd1
+ _12773_/X sky130_fd_sc_hd__a221o_1
XFILLER_187_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17300_ _17298_/Y _17299_/X _17210_/A vssd1 vssd1 vccd1 vccd1 _19450_/D sky130_fd_sc_hd__a21oi_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _17714_/A0 _18362_/Q _14517_/S vssd1 vssd1 vccd1 vccd1 _18362_/D sky130_fd_sc_hd__mux2_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _17533_/A _11724_/B vssd1 vssd1 vccd1 vccd1 _11724_/Y sky130_fd_sc_hd__nor2_4
X_18280_ _18734_/CLK _18280_/D vssd1 vssd1 vccd1 vccd1 _18280_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _19441_/Q _15124_/B _17211_/A _15491_/X vssd1 vssd1 vccd1 vccd1 _15492_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17231_/A _17231_/B vssd1 vssd1 vccd1 vccd1 _19427_/D sky130_fd_sc_hd__nor2_1
XFILLER_159_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14443_ _18582_/Q _14452_/B vssd1 vssd1 vccd1 vccd1 _18295_/D sky130_fd_sc_hd__and2_1
X_11655_ _11820_/A _11810_/A vssd1 vssd1 vccd1 vccd1 _11801_/A sky130_fd_sc_hd__nand2_8
XFILLER_230_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_88_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18627_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10606_ _10085_/A _10605_/X _11143_/A1 vssd1 vssd1 vccd1 vccd1 _10606_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17162_ _17231_/A _17162_/B vssd1 vssd1 vccd1 vccd1 _19405_/D sky130_fd_sc_hd__nor2_1
X_11586_ _18470_/Q _10838_/B _11585_/X vssd1 vssd1 vccd1 vccd1 _11586_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14374_ _18226_/Q _16548_/A0 _14377_/S vssd1 vssd1 vccd1 vccd1 _18226_/D sky130_fd_sc_hd__mux2_1
XFILLER_196_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16113_ _18759_/Q _16137_/B vssd1 vssd1 vccd1 vccd1 _16113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10537_ _11312_/A1 _19219_/Q _19187_/Q _09108_/B _11584_/C1 vssd1 vssd1 vccd1 vccd1
+ _10537_/X sky130_fd_sc_hd__a221o_1
X_13325_ _18113_/Q _13326_/B vssd1 vssd1 vccd1 vccd1 _13397_/C sky130_fd_sc_hd__and2_2
Xclkbuf_leaf_17_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19163_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_183_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17093_ _19380_/Q _17115_/B vssd1 vssd1 vccd1 vccd1 _17093_/X sky130_fd_sc_hd__or2_1
XFILLER_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16044_ _16046_/A _16044_/B vssd1 vssd1 vccd1 vccd1 _18733_/D sky130_fd_sc_hd__and2_1
X_10468_ _10466_/X _10467_/X _10618_/S vssd1 vssd1 vccd1 vccd1 _10468_/X sky130_fd_sc_hd__mux2_1
X_13256_ _09193_/X _12762_/Y _13255_/X _13256_/B1 _17930_/Q vssd1 vssd1 vccd1 vccd1
+ _13257_/B sky130_fd_sc_hd__a32o_1
XFILLER_170_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12207_ _17866_/Q _12208_/C _17867_/Q vssd1 vssd1 vccd1 vccd1 _12209_/B sky130_fd_sc_hd__a21oi_1
XFILLER_142_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13187_ _13257_/A _13187_/B vssd1 vssd1 vccd1 vccd1 _17928_/D sky130_fd_sc_hd__and2_1
XFILLER_269_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10399_ _10399_/A _10399_/B vssd1 vssd1 vccd1 vccd1 _10399_/Y sky130_fd_sc_hd__nand2_2
XFILLER_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12138_ _17841_/Q _12138_/B vssd1 vssd1 vccd1 vccd1 _12144_/C sky130_fd_sc_hd__and2_2
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17995_ _18543_/CLK _17995_/D vssd1 vssd1 vccd1 vccd1 _17995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16946_ _16848_/S _17945_/Q _16945_/X vssd1 vssd1 vccd1 vccd1 _17196_/B sky130_fd_sc_hd__o21a_4
X_12069_ _17812_/Q _12087_/B vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__or2_1
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16877_ _18750_/Q _12276_/A _16877_/B1 input245/X _12483_/A vssd1 vssd1 vccd1 vccd1
+ _16877_/X sky130_fd_sc_hd__a221o_1
XFILLER_38_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18616_ _19146_/CLK _18616_/D vssd1 vssd1 vccd1 vccd1 _18616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_252_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _18620_/Q _17718_/A0 _15833_/S vssd1 vssd1 vccd1 vccd1 _18620_/D sky130_fd_sc_hd__mux2_1
X_19596_ _19596_/CLK _19596_/D vssd1 vssd1 vccd1 vccd1 _19596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18547_ _19601_/CLK _18547_/D vssd1 vssd1 vccd1 vccd1 _18547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15759_ _19485_/Q _15758_/X _15781_/S vssd1 vssd1 vccd1 vccd1 _15759_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09280_ _09643_/A _11808_/A _09279_/Y _09946_/B1 vssd1 vssd1 vccd1 vccd1 _12600_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_205_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18478_ _19320_/CLK _18478_/D vssd1 vssd1 vccd1 vccd1 _18478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17429_ _19497_/Q _17453_/B _17427_/X _17428_/Y _17338_/A vssd1 vssd1 vccd1 vccd1
+ _19497_/D sky130_fd_sc_hd__o221a_1
XFILLER_220_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08995_ _17920_/Q _08995_/B vssd1 vssd1 vccd1 vccd1 _09245_/C sky130_fd_sc_hd__nor2_2
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09616_ _10315_/S _09615_/X _10260_/B1 vssd1 vssd1 vccd1 vccd1 _09616_/X sky130_fd_sc_hd__o21a_1
XFILLER_284_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09547_ _12471_/A0 _09545_/X _09546_/X vssd1 vssd1 vccd1 vccd1 _09547_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09478_ _11691_/B1 _09991_/A _09477_/X _11692_/A1 _18379_/Q vssd1 vssd1 vccd1 vccd1
+ _09478_/X sky130_fd_sc_hd__o32a_1
XFILLER_54_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _08958_/X _11439_/X _11376_/B _11518_/B2 vssd1 vssd1 vccd1 vccd1 _15380_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11371_ _17965_/Q _11447_/A2 _11371_/B1 vssd1 vssd1 vccd1 vccd1 _11371_/X sky130_fd_sc_hd__a21o_1
XFILLER_192_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10322_ _18870_/Q _18902_/Q _10687_/S vssd1 vssd1 vccd1 vccd1 _10322_/X sky130_fd_sc_hd__mux2_1
X_13110_ _19431_/Q _12560_/B _13108_/X _13109_/X _12560_/A vssd1 vssd1 vccd1 vccd1
+ _13110_/X sky130_fd_sc_hd__o221a_2
XFILLER_124_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14090_ _16540_/A0 _18030_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _18030_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13041_ _12815_/A _12820_/X _13041_/S vssd1 vssd1 vccd1 vccd1 _13354_/B sky130_fd_sc_hd__mux2_1
X_10253_ _10253_/A _18807_/Q _10253_/C vssd1 vssd1 vccd1 vccd1 _10253_/X sky130_fd_sc_hd__and3_1
XFILLER_152_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10184_ _10182_/X _10183_/X _10335_/S vssd1 vssd1 vccd1 vccd1 _10184_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1202 _12755_/X vssd1 vssd1 vccd1 vccd1 _13230_/A1 sky130_fd_sc_hd__buf_2
Xfanout1213 _12729_/B vssd1 vssd1 vccd1 vccd1 _13911_/A sky130_fd_sc_hd__buf_6
XFILLER_182_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1224 _15382_/B2 vssd1 vssd1 vccd1 vccd1 _15429_/A2 sky130_fd_sc_hd__buf_4
X_16800_ _16803_/A _16800_/B _16802_/B vssd1 vssd1 vccd1 vccd1 _19288_/D sky130_fd_sc_hd__nor3_1
Xfanout1235 _12265_/Y vssd1 vssd1 vccd1 vccd1 _13227_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout1246 _08944_/Y vssd1 vssd1 vccd1 vccd1 _08947_/B sky130_fd_sc_hd__buf_6
X_17780_ _19211_/CLK _17780_/D vssd1 vssd1 vccd1 vccd1 _17780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_135_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19363_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14992_ _14992_/A1 _13928_/X _14683_/X _18656_/Q vssd1 vssd1 vccd1 vccd1 _14992_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1257 _11441_/B vssd1 vssd1 vccd1 vccd1 _11490_/B sky130_fd_sc_hd__clkbuf_8
Xfanout1268 _14591_/A2 vssd1 vssd1 vccd1 vccd1 _14559_/A2 sky130_fd_sc_hd__buf_4
XFILLER_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1279 _11712_/X vssd1 vssd1 vccd1 vccd1 _11715_/B sky130_fd_sc_hd__buf_6
XFILLER_247_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16731_ _19263_/Q _16734_/C _16737_/A vssd1 vssd1 vccd1 vccd1 _16731_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13943_ _19263_/Q _13943_/A2 _13943_/B1 _19295_/Q vssd1 vssd1 vccd1 vccd1 _13943_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19450_ _19450_/CLK _19450_/D vssd1 vssd1 vccd1 vccd1 _19450_/Q sky130_fd_sc_hd__dfxtp_1
X_16662_ _16768_/A _16662_/B _16667_/C vssd1 vssd1 vccd1 vccd1 _19242_/D sky130_fd_sc_hd__nor3_1
XFILLER_235_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13874_ _13874_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _13874_/X sky130_fd_sc_hd__and2_1
XFILLER_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18401_ _19466_/CLK _18401_/D vssd1 vssd1 vccd1 vccd1 _18401_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_223_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15613_ _19478_/Q _15612_/Y _15716_/S vssd1 vssd1 vccd1 vccd1 _15613_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12825_ _12822_/Y _12824_/Y _12933_/A vssd1 vssd1 vccd1 vccd1 _12826_/A sky130_fd_sc_hd__mux2_1
X_19381_ _19477_/CLK _19381_/D vssd1 vssd1 vccd1 vccd1 _19381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16593_ _16593_/A0 _19196_/Q _16622_/S vssd1 vssd1 vccd1 vccd1 _19196_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18332_ _19611_/CLK _18332_/D vssd1 vssd1 vccd1 vccd1 _18332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ _15544_/A _15544_/B vssd1 vssd1 vccd1 vccd1 _15544_/X sky130_fd_sc_hd__xor2_1
XFILLER_188_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12756_/A _12756_/B vssd1 vssd1 vccd1 vccd1 _12756_/Y sky130_fd_sc_hd__nand2_8
XFILLER_203_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18263_ _19608_/CLK _18263_/D vssd1 vssd1 vccd1 vccd1 _18263_/Q sky130_fd_sc_hd__dfxtp_1
X_11707_ _18531_/Q _18530_/Q vssd1 vssd1 vccd1 vccd1 _11707_/X sky130_fd_sc_hd__or2_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15475_ _19472_/Q _15474_/Y _15498_/S vssd1 vssd1 vccd1 vccd1 _15475_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12687_ _12601_/B _12658_/B _13911_/A vssd1 vssd1 vccd1 vccd1 _12687_/X sky130_fd_sc_hd__mux2_2
X_17214_ _17214_/A _17214_/B vssd1 vssd1 vccd1 vccd1 _17214_/Y sky130_fd_sc_hd__nand2_1
X_14426_ _18565_/Q _16046_/A vssd1 vssd1 vccd1 vccd1 _18278_/D sky130_fd_sc_hd__and2_1
X_18194_ _19225_/CLK _18194_/D vssd1 vssd1 vccd1 vccd1 _18194_/Q sky130_fd_sc_hd__dfxtp_1
X_11638_ _11638_/A _13812_/A vssd1 vssd1 vccd1 vccd1 _13810_/A sky130_fd_sc_hd__xor2_4
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17145_ _17151_/A _17575_/A vssd1 vssd1 vccd1 vccd1 _17433_/A sky130_fd_sc_hd__nand2_1
X_14357_ _18209_/Q _17664_/A0 _14377_/S vssd1 vssd1 vccd1 vccd1 _18209_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _18657_/Q _18079_/Q _19098_/Q _19002_/Q _11226_/S _11569_/S1 vssd1 vssd1
+ vccd1 vccd1 _11569_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13308_ _13757_/A _13998_/B _13295_/Y vssd1 vssd1 vccd1 vccd1 _13321_/B sky130_fd_sc_hd__o21a_1
XFILLER_128_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17076_ _17581_/A _17114_/A2 _17075_/X _17346_/A vssd1 vssd1 vccd1 vccd1 _19371_/D
+ sky130_fd_sc_hd__o211a_1
X_14288_ _17706_/A0 _18147_/Q _14305_/S vssd1 vssd1 vccd1 vccd1 _18147_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16027_ _16020_/A _16056_/B _18728_/Q vssd1 vssd1 vccd1 vccd1 _16027_/X sky130_fd_sc_hd__a21o_1
X_13239_ _17833_/Q _13942_/A2 _13942_/B1 _17865_/Q vssd1 vssd1 vccd1 vccd1 _13239_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17978_ _18627_/CLK _17978_/D vssd1 vssd1 vccd1 vccd1 _17978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16929_ _18763_/Q _16969_/A2 _16969_/B1 input228/X _16969_/C1 vssd1 vssd1 vccd1 vccd1
+ _16929_/X sky130_fd_sc_hd__a221o_4
Xfanout1780 _17907_/Q vssd1 vssd1 vccd1 vccd1 _12320_/B sky130_fd_sc_hd__buf_12
XFILLER_284_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1791 _12389_/A1 vssd1 vssd1 vccd1 vccd1 _10742_/A1 sky130_fd_sc_hd__buf_12
XFILLER_266_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19648_ _19648_/CLK _19648_/D vssd1 vssd1 vccd1 vccd1 _19648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09401_ _09401_/A _09401_/B _09401_/C vssd1 vssd1 vccd1 vccd1 _13154_/S sky130_fd_sc_hd__or3_4
XFILLER_198_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19579_ _19611_/CLK _19579_/D vssd1 vssd1 vccd1 vccd1 _19579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09332_ _09049_/Y _09331_/Y _09328_/X _09987_/A vssd1 vssd1 vccd1 vccd1 _09332_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09263_ _09272_/A1 _18603_/Q _18174_/Q _09252_/S vssd1 vssd1 vccd1 vccd1 _09263_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09194_ _10219_/A1 _19205_/Q _19173_/Q _10128_/B _10293_/B1 vssd1 vssd1 vccd1 vccd1
+ _09194_/X sky130_fd_sc_hd__a221o_1
XFILLER_194_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08978_ _18247_/Q _18822_/Q _18450_/Q _18351_/Q _09306_/S _11510_/S1 vssd1 vssd1
+ vccd1 vccd1 _08979_/B sky130_fd_sc_hd__mux4_1
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10940_ _18862_/Q _18894_/Q _10940_/S vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10871_ _10532_/A _14510_/A0 _11800_/B vssd1 vssd1 vccd1 vccd1 _10871_/X sky130_fd_sc_hd__o21a_1
XFILLER_204_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _12610_/A _12610_/B vssd1 vssd1 vccd1 vccd1 _13033_/B sky130_fd_sc_hd__nand2_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _19348_/Q _13883_/A2 _13883_/B1 _19476_/Q _13883_/C1 vssd1 vssd1 vccd1 vccd1
+ _13590_/X sky130_fd_sc_hd__a221o_1
XFILLER_243_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _12545_/A _13167_/A vssd1 vssd1 vccd1 vccd1 _12541_/Y sky130_fd_sc_hd__nor2_1
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _15304_/A1 _13162_/B _15285_/A3 _15259_/Y vssd1 vssd1 vccd1 vccd1 _15260_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_200_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12472_ _12851_/B _12528_/C vssd1 vssd1 vccd1 vccd1 _12514_/A sky130_fd_sc_hd__nor2_4
XFILLER_61_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14211_ _18277_/Q _14252_/B _14210_/Y _16046_/A vssd1 vssd1 vccd1 vccd1 _18103_/D
+ sky130_fd_sc_hd__o211a_1
X_11423_ _09374_/S _11422_/X _11501_/B1 vssd1 vssd1 vccd1 vccd1 _11423_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15191_ _17382_/A _15190_/X _15424_/C1 vssd1 vssd1 vccd1 vccd1 _15191_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 _18287_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11354_ _11352_/X _11353_/X _11361_/S vssd1 vssd1 vccd1 vccd1 _11354_/X sky130_fd_sc_hd__mux2_1
X_14142_ _14142_/A _14142_/B _14142_/C _14141_/Y vssd1 vssd1 vccd1 vccd1 _14143_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_4_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10305_ _18129_/Q _13843_/A _13904_/A vssd1 vssd1 vccd1 vccd1 _12658_/B sky130_fd_sc_hd__mux2_4
X_18950_ _19079_/CLK _18950_/D vssd1 vssd1 vccd1 vccd1 _18950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14073_ _17690_/A0 _18015_/Q _14073_/S vssd1 vssd1 vccd1 vccd1 _18015_/D sky130_fd_sc_hd__mux2_1
X_11285_ _11283_/X _11284_/X _11285_/S vssd1 vssd1 vccd1 vccd1 _11285_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13024_ _13303_/B2 _13009_/X _13012_/X _13023_/X vssd1 vssd1 vccd1 vccd1 _13024_/X
+ sky130_fd_sc_hd__a22o_4
X_10236_ _17980_/Q _11447_/A2 _11371_/B1 vssd1 vssd1 vccd1 vccd1 _10236_/X sky130_fd_sc_hd__a21o_1
X_17901_ _17901_/CLK _17901_/D vssd1 vssd1 vccd1 vccd1 _17901_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_239_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18881_ _18881_/CLK _18881_/D vssd1 vssd1 vccd1 vccd1 _18881_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1010 _16459_/X vssd1 vssd1 vccd1 vccd1 _16488_/S sky130_fd_sc_hd__buf_8
XFILLER_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1021 _14973_/A1 vssd1 vssd1 vccd1 vccd1 _14992_/A1 sky130_fd_sc_hd__buf_6
X_17832_ _17865_/CLK _17832_/D vssd1 vssd1 vccd1 vccd1 _17832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_266_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10167_ _19647_/Q _18936_/Q _10168_/S vssd1 vssd1 vccd1 vccd1 _10167_/X sky130_fd_sc_hd__mux2_1
Xfanout1032 _16465_/A0 vssd1 vssd1 vccd1 vccd1 _16597_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout1043 _15081_/A vssd1 vssd1 vccd1 vccd1 _11816_/A sky130_fd_sc_hd__buf_12
XFILLER_255_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1054 _17559_/X vssd1 vssd1 vccd1 vccd1 _17603_/B1 sky130_fd_sc_hd__buf_6
Xfanout1065 _13486_/A1 vssd1 vssd1 vccd1 vccd1 _13312_/A sky130_fd_sc_hd__buf_4
XFILLER_120_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17763_ _19608_/CLK _17763_/D vssd1 vssd1 vccd1 vccd1 _17763_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1076 _17659_/A0 vssd1 vssd1 vccd1 vccd1 _17692_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_282_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10098_ _18266_/Q _18841_/Q _10099_/S vssd1 vssd1 vccd1 vccd1 _10098_/X sky130_fd_sc_hd__mux2_1
X_14975_ _18129_/Q _14671_/X _14934_/X _14974_/X vssd1 vssd1 vccd1 vccd1 _14975_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout1087 _09825_/X vssd1 vssd1 vccd1 vccd1 _16462_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1098 _17516_/C1 vssd1 vssd1 vccd1 vccd1 _08883_/A sky130_fd_sc_hd__buf_6
XFILLER_281_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16714_ _16808_/A _16714_/B _16715_/B vssd1 vssd1 vccd1 vccd1 _19257_/D sky130_fd_sc_hd__nor3_1
X_19502_ _19502_/CLK _19502_/D vssd1 vssd1 vccd1 vccd1 _19502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13926_ _19326_/Q _13165_/C _12584_/B _13181_/Y _13925_/X vssd1 vssd1 vccd1 vccd1
+ _13926_/X sky130_fd_sc_hd__o32a_2
XFILLER_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17694_ _17694_/A0 _19620_/Q _17723_/S vssd1 vssd1 vccd1 vccd1 _19620_/D sky130_fd_sc_hd__mux2_1
XFILLER_281_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19433_ _19433_/CLK _19433_/D vssd1 vssd1 vccd1 vccd1 _19433_/Q sky130_fd_sc_hd__dfxtp_1
X_16645_ _19237_/Q _16641_/B _16644_/Y vssd1 vssd1 vccd1 vccd1 _19237_/D sky130_fd_sc_hd__o21a_1
XFILLER_235_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13857_ _13637_/A _14030_/B _13843_/Y vssd1 vssd1 vccd1 vccd1 _13857_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19364_ _19522_/CLK _19364_/D vssd1 vssd1 vccd1 vccd1 _19364_/Q sky130_fd_sc_hd__dfxtp_1
X_12808_ _12799_/X _12807_/X _13354_/A vssd1 vssd1 vccd1 vccd1 _12808_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16576_ _17676_/A0 _19180_/Q _16585_/S vssd1 vssd1 vccd1 vccd1 _19180_/D sky130_fd_sc_hd__mux2_1
X_13788_ _14026_/B vssd1 vssd1 vccd1 vccd1 _13788_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18315_ _19126_/CLK _18315_/D vssd1 vssd1 vccd1 vccd1 _18315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15527_ _15526_/B _13576_/Y _15133_/B _15526_/Y vssd1 vssd1 vccd1 vccd1 _15527_/X
+ sky130_fd_sc_hd__a31o_1
X_19295_ _19295_/CLK _19295_/D vssd1 vssd1 vccd1 vccd1 _19295_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_32_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19634_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12739_ _12702_/Y _12738_/Y _12739_/S vssd1 vssd1 vccd1 vccd1 _12739_/X sky130_fd_sc_hd__mux2_2
XFILLER_188_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18246_ _19126_/CLK _18246_/D vssd1 vssd1 vccd1 vccd1 _18246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15458_ _15364_/A _15364_/B _15457_/A vssd1 vssd1 vccd1 vccd1 _15458_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14409_ _17716_/A0 _18260_/Q _14416_/S vssd1 vssd1 vccd1 vccd1 _18260_/D sky130_fd_sc_hd__mux2_1
X_18177_ _19630_/CLK _18177_/D vssd1 vssd1 vccd1 vccd1 _18177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ _18574_/Q _15388_/C _18575_/Q vssd1 vssd1 vccd1 vccd1 _15390_/B sky130_fd_sc_hd__a21oi_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17128_ _19394_/Q _17120_/Y _17127_/X vssd1 vssd1 vccd1 vccd1 _19394_/D sky130_fd_sc_hd__o21ba_1
XFILLER_237_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09950_ _11497_/A1 _19196_/Q _19164_/Q _09973_/S _10144_/B1 vssd1 vssd1 vccd1 vccd1
+ _09950_/X sky130_fd_sc_hd__a221o_1
X_17059_ _17565_/B _17113_/B vssd1 vssd1 vccd1 vccd1 _17059_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08901_ _08901_/A _12023_/A vssd1 vssd1 vccd1 vccd1 _08901_/Y sky130_fd_sc_hd__nor2_2
XFILLER_170_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _08901_/A _19556_/Q _10054_/S _19588_/Q _10033_/S vssd1 vssd1 vccd1 vccd1
+ _09881_/X sky130_fd_sc_hd__o221a_1
XFILLER_258_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08832_ _18124_/Q vssd1 vssd1 vccd1 vccd1 _14252_/A sky130_fd_sc_hd__inv_2
XFILLER_285_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09315_ _09317_/B vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__inv_2
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09246_ _09049_/Y _09903_/B _09241_/Y _09987_/A vssd1 vssd1 vccd1 vccd1 _09246_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_193_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09177_ _18246_/Q _18821_/Q _18449_/Q _18350_/Q _09344_/S _08843_/A vssd1 vssd1 vccd1
+ vccd1 _09177_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11070_ _18643_/Q _18065_/Q _11070_/S vssd1 vssd1 vccd1 vccd1 _11070_/X sky130_fd_sc_hd__mux2_1
XFILLER_277_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput102 dout0[63] vssd1 vssd1 vccd1 vccd1 input102/X sky130_fd_sc_hd__clkbuf_2
X_10021_ _09095_/A _10017_/X _10020_/X vssd1 vssd1 vccd1 vccd1 _10021_/X sky130_fd_sc_hd__a21o_1
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput113 dout1[15] vssd1 vssd1 vccd1 vccd1 input113/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput124 dout1[25] vssd1 vssd1 vccd1 vccd1 input124/X sky130_fd_sc_hd__clkbuf_2
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput135 dout1[35] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_hd__buf_2
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput146 dout1[45] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_hd__clkbuf_2
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput157 dout1[55] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_hd__buf_2
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 dout1[7] vssd1 vssd1 vccd1 vccd1 input168/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 irq[2] vssd1 vssd1 vccd1 vccd1 input179/X sky130_fd_sc_hd__clkbuf_4
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _14992_/A1 _13118_/Y _14973_/B1 _18633_/Q _14741_/B vssd1 vssd1 vccd1 vccd1
+ _14760_/X sky130_fd_sc_hd__a221o_2
XFILLER_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11972_ _18737_/Q _18736_/Q _18735_/Q _11972_/D vssd1 vssd1 vccd1 vccd1 _11972_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _13711_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13711_/Y sky130_fd_sc_hd__nor2_1
XFILLER_189_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _18035_/Q _18003_/Q _11309_/S vssd1 vssd1 vccd1 vccd1 _10923_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _18101_/Q _14801_/B _14684_/X _14690_/Y vssd1 vssd1 vccd1 vccd1 _14691_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_244_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16430_ _19038_/Q _17695_/A0 _16453_/S vssd1 vssd1 vccd1 vccd1 _19038_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13642_ _18122_/Q _13642_/B vssd1 vssd1 vccd1 vccd1 _13643_/B sky130_fd_sc_hd__nor2_1
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10854_ _10852_/X _10853_/X _11577_/S vssd1 vssd1 vccd1 vccd1 _10854_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16461_/A0 _18972_/Q _16388_/S vssd1 vssd1 vccd1 vccd1 _18972_/D sky130_fd_sc_hd__mux2_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13573_ _13566_/Y _13569_/Y _13571_/Y _13572_/X vssd1 vssd1 vccd1 vccd1 _13573_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ _10785_/A _10785_/B vssd1 vssd1 vccd1 vccd1 _10785_/X sky130_fd_sc_hd__or2_1
X_18100_ _18713_/CLK _18100_/D vssd1 vssd1 vccd1 vccd1 _18100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15365_/C _15312_/B vssd1 vssd1 vccd1 vccd1 _15313_/B sky130_fd_sc_hd__nand2_1
X_19080_ _19565_/CLK _19080_/D vssd1 vssd1 vccd1 vccd1 _19080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12524_ _12577_/B _12768_/B vssd1 vssd1 vccd1 vccd1 _12524_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _16292_/A0 _18906_/Q _16292_/S vssd1 vssd1 vccd1 vccd1 _18906_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18031_ _19601_/CLK _18031_/D vssd1 vssd1 vccd1 vccd1 _18031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15243_ _15243_/A _15243_/B vssd1 vssd1 vccd1 vccd1 _15263_/D sky130_fd_sc_hd__xor2_4
X_12455_ _12455_/A _12587_/B vssd1 vssd1 vccd1 vccd1 _12455_/Y sky130_fd_sc_hd__nand2_2
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11406_ _11400_/X _11402_/X _11405_/X _11406_/B2 _09350_/S vssd1 vssd1 vccd1 vccd1
+ _11406_/X sky130_fd_sc_hd__o221a_2
XFILLER_172_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15174_ _15259_/B _12982_/B _15285_/A3 _15173_/Y vssd1 vssd1 vccd1 vccd1 _15174_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12386_ _17903_/Q _12408_/B _12385_/X _13981_/C1 vssd1 vssd1 vccd1 vccd1 _17903_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ _16476_/A0 _18064_/Q _14131_/S vssd1 vssd1 vccd1 vccd1 _18064_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11337_ _18115_/Q _11337_/B vssd1 vssd1 vccd1 vccd1 _11337_/X sky130_fd_sc_hd__or2_2
XFILLER_67_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_150_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19533_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18933_ _19644_/CLK _18933_/D vssd1 vssd1 vccd1 vccd1 _18933_/Q sky130_fd_sc_hd__dfxtp_1
X_14056_ _16540_/A0 _17998_/Q _14073_/S vssd1 vssd1 vccd1 vccd1 _17998_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ _11277_/A1 _19210_/Q _19178_/Q _11284_/B2 vssd1 vssd1 vccd1 vccd1 _11268_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13007_ _14487_/A _13007_/B vssd1 vssd1 vccd1 vccd1 _17924_/D sky130_fd_sc_hd__nor2_1
XFILLER_122_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10219_ _10219_/A1 _18162_/Q _18808_/Q _10215_/S vssd1 vssd1 vccd1 vccd1 _10219_/X
+ sky130_fd_sc_hd__a22o_1
X_11199_ _18859_/Q _18891_/Q _19051_/Q _19019_/Q _10717_/S _11199_/S1 vssd1 vssd1
+ vccd1 vccd1 _11199_/X sky130_fd_sc_hd__mux4_1
X_18864_ _19607_/CLK _18864_/D vssd1 vssd1 vccd1 vccd1 _18864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_282_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17815_ _19492_/CLK _17815_/D vssd1 vssd1 vccd1 vccd1 _17815_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18795_ _19211_/CLK _18795_/D vssd1 vssd1 vccd1 vccd1 _18795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17746_ _18646_/Q vssd1 vssd1 vccd1 vccd1 _18646_/D sky130_fd_sc_hd__clkbuf_2
X_14958_ _14958_/A vssd1 vssd1 vccd1 vccd1 _14958_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_242_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13909_ _13958_/B _14152_/C _13909_/B1 vssd1 vssd1 vccd1 vccd1 _13909_/Y sky130_fd_sc_hd__a21oi_1
X_17677_ _17677_/A0 _19604_/Q _17689_/S vssd1 vssd1 vccd1 vccd1 _19604_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14889_ _14885_/X _14888_/X _14889_/B1 vssd1 vssd1 vccd1 vccd1 _14889_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16628_ _19650_/Q _08991_/A _17887_/Q _17724_/B _12460_/A vssd1 vssd1 vccd1 vccd1
+ _16628_/X sky130_fd_sc_hd__a41o_1
X_19416_ _19482_/CLK _19416_/D vssd1 vssd1 vccd1 vccd1 _19416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19347_ _19542_/CLK _19347_/D vssd1 vssd1 vccd1 vccd1 _19347_/Q sky130_fd_sc_hd__dfxtp_1
X_16559_ _16592_/A0 _19163_/Q _16590_/S vssd1 vssd1 vccd1 vccd1 _19163_/D sky130_fd_sc_hd__mux2_1
X_09100_ _14350_/A _09857_/A1 _09106_/B _16392_/C _09094_/Y vssd1 vssd1 vccd1 vccd1
+ _09102_/C sky130_fd_sc_hd__a221o_1
X_19278_ _19280_/CLK _19278_/D vssd1 vssd1 vccd1 vccd1 _19278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09031_ _11556_/A _08996_/B _09031_/S vssd1 vssd1 vccd1 vccd1 _09032_/B sky130_fd_sc_hd__mux2_1
X_18229_ _19620_/CLK _18229_/D vssd1 vssd1 vccd1 vccd1 _18229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09933_ _19036_/Q _19004_/Q _11472_/C vssd1 vssd1 vccd1 vccd1 _09933_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout803 _16165_/S vssd1 vssd1 vccd1 vccd1 _16189_/S sky130_fd_sc_hd__buf_12
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout814 _14351_/Y vssd1 vssd1 vccd1 vccd1 _14377_/S sky130_fd_sc_hd__clkbuf_16
Xfanout825 _12762_/Y vssd1 vssd1 vccd1 vccd1 _13292_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_259_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout836 _16543_/A0 vssd1 vssd1 vccd1 vccd1 _16609_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout847 _14510_/A0 vssd1 vssd1 vccd1 vccd1 _16314_/A0 sky130_fd_sc_hd__clkbuf_4
X_09864_ _09862_/X _09863_/Y _09141_/A vssd1 vssd1 vccd1 vccd1 _12602_/A sky130_fd_sc_hd__a21oi_4
Xfanout858 _10713_/A2 vssd1 vssd1 vccd1 vccd1 _17681_/A0 sky130_fd_sc_hd__clkbuf_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout869 _16455_/A1 vssd1 vssd1 vccd1 vccd1 _17720_/A0 sky130_fd_sc_hd__clkbuf_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08815_ _19650_/Q vssd1 vssd1 vccd1 vccd1 _17724_/A sky130_fd_sc_hd__inv_6
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09795_ _09783_/X _09794_/X _11607_/S vssd1 vssd1 vccd1 vccd1 _09795_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_207 _18778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 _17914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _18387_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10570_ _18040_/Q _18008_/Q _10645_/S vssd1 vssd1 vccd1 vccd1 _10570_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09229_ _12599_/A _09229_/B vssd1 vssd1 vccd1 vccd1 _09230_/B sky130_fd_sc_hd__nand2_2
XFILLER_194_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ _17878_/Q _17879_/Q _12240_/C vssd1 vssd1 vccd1 vccd1 _12242_/B sky130_fd_sc_hd__and3_1
XFILLER_181_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12171_ _16811_/A _12176_/C vssd1 vssd1 vccd1 vccd1 _12171_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11122_ _11112_/A _11121_/X _11608_/C1 vssd1 vssd1 vccd1 vccd1 _11122_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15930_ _18685_/Q _15948_/A2 _15923_/C _15929_/X _15945_/C1 vssd1 vssd1 vccd1 vccd1
+ _15930_/X sky130_fd_sc_hd__a221o_1
X_11053_ _11053_/A _11053_/B _11053_/C vssd1 vssd1 vccd1 vccd1 _11053_/X sky130_fd_sc_hd__or3_1
XFILLER_277_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10004_ _10004_/A1 _09999_/X _10000_/X _10003_/X _11570_/B1 vssd1 vssd1 vccd1 vccd1
+ _10009_/B sky130_fd_sc_hd__o311a_1
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15861_ _18662_/Q _15853_/Y _15906_/B1 vssd1 vssd1 vccd1 vccd1 _15861_/X sky130_fd_sc_hd__a21o_1
XFILLER_236_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17600_ _19541_/Q _17624_/A2 _17599_/X _17356_/A vssd1 vssd1 vccd1 vccd1 _19541_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _14964_/B1 _14810_/X _14811_/X _14771_/X vssd1 vssd1 vccd1 vccd1 _14812_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _19521_/CLK _18580_/D vssd1 vssd1 vccd1 vccd1 _18580_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_76_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _15793_/A2 _15790_/X _15791_/Y _15623_/A vssd1 vssd1 vccd1 vccd1 _15792_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_224_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _17531_/A _17531_/B vssd1 vssd1 vccd1 vccd1 _17531_/Y sky130_fd_sc_hd__nor2_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _14741_/Y _14742_/X _14964_/B1 vssd1 vssd1 vccd1 vccd1 _14743_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11955_ _19228_/Q _11959_/A2 _14343_/C _11959_/B2 vssd1 vssd1 vccd1 vccd1 _11955_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10906_ _10908_/B vssd1 vssd1 vccd1 vccd1 _12641_/B sky130_fd_sc_hd__inv_2
XFILLER_60_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17462_ _17462_/A _17462_/B vssd1 vssd1 vccd1 vccd1 _17462_/Y sky130_fd_sc_hd__nand2_1
XFILLER_264_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14674_ _17790_/Q _14911_/B vssd1 vssd1 vccd1 vccd1 _14674_/X sky130_fd_sc_hd__or2_1
XFILLER_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11886_ _11899_/A _11886_/B _11886_/C vssd1 vssd1 vccd1 vccd1 _11886_/X sky130_fd_sc_hd__and3_4
XFILLER_205_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19201_ _19201_/CLK _19201_/D vssd1 vssd1 vccd1 vccd1 _19201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16413_ _16611_/A0 _19022_/Q _16420_/S vssd1 vssd1 vccd1 vccd1 _19022_/D sky130_fd_sc_hd__mux2_1
X_13625_ _19253_/Q _13625_/A2 _13625_/B1 _19285_/Q vssd1 vssd1 vccd1 vccd1 _13625_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_177_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10837_ _17940_/Q _11451_/A2 _10836_/X _08947_/B vssd1 vssd1 vccd1 vccd1 _10837_/X
+ sky130_fd_sc_hd__o22a_4
X_17393_ _18101_/Q _17546_/A2 _17392_/X vssd1 vssd1 vccd1 vccd1 _17393_/X sky130_fd_sc_hd__o21a_2
XFILLER_186_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19132_ _19587_/CLK _19132_/D vssd1 vssd1 vccd1 vccd1 _19132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16344_ _18956_/Q _16543_/A0 _16358_/S vssd1 vssd1 vccd1 vccd1 _18956_/D sky130_fd_sc_hd__mux2_1
X_13556_ _19443_/Q _13949_/A2 _13554_/X _13555_/X _13949_/C1 vssd1 vssd1 vccd1 vccd1
+ _13556_/X sky130_fd_sc_hd__o221a_1
XFILLER_201_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10768_ _18257_/Q _18832_/Q _11576_/S vssd1 vssd1 vccd1 vccd1 _10768_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19063_ _19625_/CLK _19063_/D vssd1 vssd1 vccd1 vccd1 _19063_/Q sky130_fd_sc_hd__dfxtp_1
X_12507_ _12507_/A _12528_/C vssd1 vssd1 vccd1 vccd1 _12576_/A sky130_fd_sc_hd__nand2_4
XFILLER_157_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16275_ _16606_/A0 _18889_/Q _16292_/S vssd1 vssd1 vccd1 vccd1 _18889_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13487_ _14155_/B _12756_/Y _13487_/S vssd1 vssd1 vccd1 vccd1 _13487_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10699_ _11250_/A1 _19576_/Q _10687_/S _19608_/Q vssd1 vssd1 vccd1 vccd1 _10699_/X
+ sky130_fd_sc_hd__o22a_1
X_18014_ _19648_/CLK _18014_/D vssd1 vssd1 vccd1 vccd1 _18014_/Q sky130_fd_sc_hd__dfxtp_1
X_15226_ _15270_/C _15226_/B vssd1 vssd1 vccd1 vccd1 _15226_/X sky130_fd_sc_hd__or2_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12438_ _17894_/Q _12438_/B vssd1 vssd1 vccd1 vccd1 _12443_/C sky130_fd_sc_hd__or2_2
XFILLER_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput406 _11928_/X vssd1 vssd1 vccd1 vccd1 din0[8] sky130_fd_sc_hd__buf_4
Xoutput417 _18487_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[16] sky130_fd_sc_hd__buf_4
XFILLER_5_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput428 _18497_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[26] sky130_fd_sc_hd__buf_4
X_15157_ _15135_/A _15135_/B _15155_/A _15155_/B vssd1 vssd1 vccd1 vccd1 _15157_/X
+ sky130_fd_sc_hd__a22o_1
X_12369_ _18383_/Q _12417_/B1 _09154_/Y _08858_/A vssd1 vssd1 vccd1 vccd1 _12370_/B
+ sky130_fd_sc_hd__a2bb2o_2
Xoutput439 _18478_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[7] sky130_fd_sc_hd__buf_4
XFILLER_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14108_ _16525_/A _16393_/A vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__nand2_8
X_15088_ _19387_/Q _15088_/B _15088_/C vssd1 vssd1 vccd1 vccd1 _15088_/X sky130_fd_sc_hd__and3_1
XFILLER_80_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18916_ _19627_/CLK _18916_/D vssd1 vssd1 vccd1 vccd1 _18916_/Q sky130_fd_sc_hd__dfxtp_1
X_14039_ _17798_/Q _14074_/C _16459_/B vssd1 vssd1 vccd1 vccd1 _16393_/A sky130_fd_sc_hd__nor3_4
XFILLER_80_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18847_ _19138_/CLK _18847_/D vssd1 vssd1 vccd1 vccd1 _18847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09580_ _18241_/Q _18816_/Q _10362_/S vssd1 vssd1 vccd1 vccd1 _09580_/X sky130_fd_sc_hd__mux2_1
XFILLER_282_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18778_ _18778_/CLK _18778_/D vssd1 vssd1 vccd1 vccd1 _18778_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_227_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17729_ _18629_/Q vssd1 vssd1 vccd1 vccd1 _18629_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_36_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09014_ _09245_/A _09031_/S vssd1 vssd1 vccd1 vccd1 _11141_/A sky130_fd_sc_hd__or2_4
XFILLER_128_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout600 _14244_/B vssd1 vssd1 vccd1 vccd1 _14260_/B sky130_fd_sc_hd__buf_4
Xfanout611 _11926_/A1 vssd1 vssd1 vccd1 vccd1 _11887_/B1 sky130_fd_sc_hd__buf_8
Xfanout1609 _15103_/Y vssd1 vssd1 vccd1 vccd1 _17461_/A2 sky130_fd_sc_hd__buf_6
X_09916_ _10262_/A1 _19555_/Q _09925_/S _19587_/Q _10337_/S1 vssd1 vssd1 vccd1 vccd1
+ _09916_/X sky130_fd_sc_hd__o221a_1
XFILLER_160_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout622 _17032_/A2 vssd1 vssd1 vccd1 vccd1 _17046_/A2 sky130_fd_sc_hd__buf_6
Xfanout633 _11818_/A vssd1 vssd1 vccd1 vccd1 _11810_/A sky130_fd_sc_hd__buf_12
Xfanout644 _17074_/A2 vssd1 vssd1 vccd1 vccd1 _17114_/A2 sky130_fd_sc_hd__buf_4
XFILLER_246_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout655 _13277_/S vssd1 vssd1 vccd1 vccd1 _13921_/S sky130_fd_sc_hd__buf_4
XFILLER_258_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout666 _12555_/Y vssd1 vssd1 vccd1 vccd1 _12570_/A sky130_fd_sc_hd__buf_6
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout677 _13246_/B1 vssd1 vssd1 vccd1 vccd1 _13950_/B1 sky130_fd_sc_hd__buf_6
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09847_ _18941_/Q _10001_/S _09853_/S _09846_/X vssd1 vssd1 vccd1 vccd1 _09847_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout688 _13654_/B1 vssd1 vssd1 vccd1 vccd1 _13948_/B1 sky130_fd_sc_hd__buf_4
XFILLER_86_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout699 _12545_/Y vssd1 vssd1 vccd1 vccd1 _13495_/B1 sky130_fd_sc_hd__buf_4
XFILLER_274_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09776_/X _09777_/Y _09946_/B1 vssd1 vssd1 vccd1 vccd1 _09816_/A sky130_fd_sc_hd__a21oi_4
XFILLER_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11740_/A vssd1 vssd1 vccd1 vccd1 _11740_/Y sky130_fd_sc_hd__inv_6
XFILLER_230_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11671_ _11671_/A _13616_/A vssd1 vssd1 vccd1 vccd1 _13622_/B sky130_fd_sc_hd__xor2_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _12626_/B _13387_/B _12596_/Y vssd1 vssd1 vccd1 vccd1 _13411_/B sky130_fd_sc_hd__o21ba_1
X_10622_ _10612_/X _10615_/X _10618_/X _10621_/X _11328_/S _11588_/B1 vssd1 vssd1
+ vccd1 vccd1 _10623_/B sky130_fd_sc_hd__mux4_2
X_14390_ _17697_/A0 _18241_/Q _14412_/S vssd1 vssd1 vccd1 vccd1 _18241_/D sky130_fd_sc_hd__mux2_1
XFILLER_169_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ input268/X _12575_/Y _13335_/X _13427_/A1 vssd1 vssd1 vccd1 vccd1 _13341_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _10633_/A _10552_/X _11563_/B1 vssd1 vssd1 vccd1 vccd1 _10553_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16060_ _18738_/Q _16063_/A _18739_/Q vssd1 vssd1 vccd1 vccd1 _16075_/B sky130_fd_sc_hd__or3b_2
XFILLER_127_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13272_ _18111_/Q _13271_/C _18112_/Q vssd1 vssd1 vccd1 vccd1 _13273_/B sky130_fd_sc_hd__a21oi_1
X_10484_ _18651_/Q _18073_/Q _19092_/Q _18996_/Q _10840_/S _10918_/C1 vssd1 vssd1
+ vccd1 vccd1 _10484_/X sky130_fd_sc_hd__mux4_1
X_15011_ _18502_/Q _15011_/A2 _15010_/Y _16803_/A vssd1 vssd1 vccd1 vccd1 _18502_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12223_ _17872_/Q _12224_/C _17873_/Q vssd1 vssd1 vccd1 vccd1 _12225_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12154_ _17847_/Q _12154_/B vssd1 vssd1 vccd1 vccd1 _12160_/C sky130_fd_sc_hd__and2_2
XFILLER_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ _18253_/Q _18828_/Q _18456_/Q _18357_/Q _11353_/B2 _11338_/S1 vssd1 vssd1
+ vccd1 vccd1 _11106_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16962_ _16970_/A1 _17949_/Q _16961_/X vssd1 vssd1 vccd1 vccd1 _17208_/B sky130_fd_sc_hd__o21a_4
XFILLER_150_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12085_ _17820_/Q _12085_/B vssd1 vssd1 vccd1 vccd1 _12085_/X sky130_fd_sc_hd__or2_1
XFILLER_249_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18701_ _18749_/CLK _18701_/D vssd1 vssd1 vccd1 vccd1 _18701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15913_ _18680_/Q _15943_/A2 _15912_/X _16764_/B1 vssd1 vssd1 vccd1 vccd1 _18680_/D
+ sky130_fd_sc_hd__o211a_1
X_11036_ _11512_/A1 _19117_/Q _19149_/Q _11426_/B2 vssd1 vssd1 vccd1 vccd1 _11036_/X
+ sky130_fd_sc_hd__a22o_1
X_16893_ _18754_/Q _16893_/A2 _16893_/B1 input218/X _12483_/A vssd1 vssd1 vccd1 vccd1
+ _16893_/X sky130_fd_sc_hd__a221o_1
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15844_ _12488_/A _15843_/A _15843_/Y _14177_/A vssd1 vssd1 vccd1 vccd1 _18660_/D
+ sky130_fd_sc_hd__o211a_1
X_18632_ _18632_/CLK _18632_/D vssd1 vssd1 vccd1 vccd1 _18632_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _19454_/Q _15793_/A2 _17208_/A _15774_/X vssd1 vssd1 vccd1 vccd1 _15775_/X
+ sky130_fd_sc_hd__o211a_1
X_18563_ _19618_/CLK _18563_/D vssd1 vssd1 vccd1 vccd1 _18563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _13349_/B _14142_/A _12986_/X vssd1 vssd1 vccd1 vccd1 _12987_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_280_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _15834_/C _14689_/Y _14854_/D vssd1 vssd1 vccd1 vccd1 _14726_/X sky130_fd_sc_hd__o21ba_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ _19514_/Q _17523_/B _17512_/X _17513_/Y _17592_/B vssd1 vssd1 vccd1 vccd1
+ _19514_/D sky130_fd_sc_hd__o221a_1
X_18494_ _19286_/CLK _18494_/D vssd1 vssd1 vccd1 vccd1 _18494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11938_ _14667_/A1 _11849_/B _11953_/A2 input224/X vssd1 vssd1 vccd1 vccd1 _11938_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17445_ _13258_/A _17445_/A2 _17445_/B1 _17801_/Q _17445_/C1 vssd1 vssd1 vccd1 vccd1
+ _17445_/X sky130_fd_sc_hd__a221o_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14657_ _17716_/A0 _18463_/Q _14664_/S vssd1 vssd1 vccd1 vccd1 _18463_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11869_ _11869_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _11869_/Y sky130_fd_sc_hd__nand2_2
XFILLER_232_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13608_ _13642_/B _13608_/B vssd1 vssd1 vccd1 vccd1 _13608_/X sky130_fd_sc_hd__or2_1
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17376_ _17376_/A _17376_/B vssd1 vssd1 vccd1 vccd1 _19485_/D sky130_fd_sc_hd__and2_1
X_14588_ _14592_/A _14588_/B vssd1 vssd1 vccd1 vccd1 _18402_/D sky130_fd_sc_hd__or2_1
XFILLER_174_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19115_ _19147_/CLK _19115_/D vssd1 vssd1 vccd1 vccd1 _19115_/Q sky130_fd_sc_hd__dfxtp_1
X_16327_ _18939_/Q _16526_/A0 _16358_/S vssd1 vssd1 vccd1 vccd1 _18939_/D sky130_fd_sc_hd__mux2_1
X_13539_ _13323_/X _13530_/X _13538_/X _13968_/B2 vssd1 vssd1 vccd1 vccd1 _13539_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_186_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19046_ _19206_/CLK _19046_/D vssd1 vssd1 vccd1 vccd1 _19046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16258_ _16622_/A0 _18873_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _18873_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15209_ _15223_/A _15206_/X _15208_/Y _15416_/A vssd1 vssd1 vccd1 vccd1 _15209_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16189_ _16619_/A0 _18806_/Q _16189_/S vssd1 vssd1 vccd1 vccd1 _18806_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09701_ _10282_/A1 _18137_/Q _18783_/Q _09704_/S _10293_/B1 vssd1 vssd1 vccd1 vccd1
+ _09701_/X sky130_fd_sc_hd__a221o_1
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09632_ _19040_/Q _19008_/Q _10320_/S vssd1 vssd1 vccd1 vccd1 _09632_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09563_ input162/X input137/X _09990_/S vssd1 vssd1 vccd1 vccd1 _09563_/X sky130_fd_sc_hd__mux2_8
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09494_ _09494_/A _18881_/Q _12024_/A vssd1 vssd1 vccd1 vccd1 _09494_/X sky130_fd_sc_hd__and3_1
XFILLER_24_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1406 fanout1407/X vssd1 vssd1 vccd1 vccd1 _09539_/S sky130_fd_sc_hd__buf_4
XFILLER_48_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1417 _11403_/S vssd1 vssd1 vccd1 vccd1 _11481_/C sky130_fd_sc_hd__clkbuf_8
Xfanout1428 _09089_/Y vssd1 vssd1 vccd1 vccd1 _09137_/S sky130_fd_sc_hd__buf_12
XFILLER_219_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1439 _09534_/S vssd1 vssd1 vccd1 vccd1 _10706_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout496 _11945_/B1 vssd1 vssd1 vccd1 vccd1 _11959_/A2 sky130_fd_sc_hd__buf_6
XFILLER_101_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12910_ _19525_/Q _19493_/Q _13372_/S vssd1 vssd1 vccd1 vccd1 _12910_/X sky130_fd_sc_hd__mux2_1
XFILLER_246_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13890_ _13860_/A _13860_/B _12658_/Y vssd1 vssd1 vccd1 vccd1 _13891_/B sky130_fd_sc_hd__a21boi_4
XFILLER_273_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ _11826_/A _13349_/B _12442_/C vssd1 vssd1 vccd1 vccd1 _12841_/X sky130_fd_sc_hd__a21o_1
XFILLER_206_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15638_/A _15556_/X _15558_/X _15580_/B _15789_/B1 vssd1 vssd1 vccd1 vccd1
+ _15560_/X sky130_fd_sc_hd__a311o_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _19523_/Q _19491_/Q _13372_/S vssd1 vssd1 vccd1 vccd1 _12772_/X sky130_fd_sc_hd__mux2_1
XFILLER_215_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _17713_/A0 _18361_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _18361_/D sky130_fd_sc_hd__mux2_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11718_/Y _11719_/X _11721_/Y vssd1 vssd1 vccd1 vccd1 _11723_/X sky130_fd_sc_hd__a21bo_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _15537_/B1 _15488_/X _15490_/Y _15751_/A vssd1 vssd1 vccd1 vccd1 _15491_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_42_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _19427_/Q _17244_/B _17229_/X vssd1 vssd1 vccd1 vccd1 _17231_/B sky130_fd_sc_hd__a21oi_1
XFILLER_230_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14442_ _18581_/Q _14442_/B vssd1 vssd1 vccd1 vccd1 _18294_/D sky130_fd_sc_hd__and2_1
XFILLER_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11654_ _11824_/A _11826_/A vssd1 vssd1 vccd1 vccd1 _11654_/Y sky130_fd_sc_hd__nor2_1
X_10605_ _09009_/X _09034_/B _09326_/A vssd1 vssd1 vccd1 vccd1 _10605_/X sky130_fd_sc_hd__a21o_1
X_17161_ _19405_/Q fanout534/X _17457_/A _17212_/B2 vssd1 vssd1 vccd1 vccd1 _17162_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14373_ _18225_/Q _17680_/A0 _14383_/S vssd1 vssd1 vccd1 vccd1 _18225_/D sky130_fd_sc_hd__mux2_1
X_11585_ _10027_/A _18371_/Q _12442_/B _11327_/S vssd1 vssd1 vccd1 vccd1 _11585_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_127_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16112_ _16078_/X _16111_/Y _12107_/A vssd1 vssd1 vccd1 vccd1 _18758_/D sky130_fd_sc_hd__a21oi_1
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13324_ _13294_/X _13321_/X _13968_/A1 _13320_/X _13968_/B2 vssd1 vssd1 vccd1 vccd1
+ _13324_/X sky130_fd_sc_hd__a32o_1
XFILLER_196_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _11252_/S _10536_/B vssd1 vssd1 vccd1 vccd1 _10536_/Y sky130_fd_sc_hd__nor2_1
X_17092_ _17178_/B _17116_/A2 _17091_/X _17356_/A vssd1 vssd1 vccd1 vccd1 _19379_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16043_ _18726_/Q _18733_/Q _16051_/S vssd1 vssd1 vccd1 vccd1 _16044_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13255_ _13255_/A _13255_/B _13234_/X vssd1 vssd1 vccd1 vccd1 _13255_/X sky130_fd_sc_hd__or3b_1
X_10467_ _18619_/Q _18190_/Q _10467_/S vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ _17866_/Q _12208_/C _12205_/Y vssd1 vssd1 vccd1 vccd1 _17866_/D sky130_fd_sc_hd__o21a_1
XFILLER_269_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_57_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19615_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_170_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13186_ _09367_/X _12762_/Y _13185_/X _13256_/B1 _17928_/Q vssd1 vssd1 vccd1 vccd1
+ _13187_/B sky130_fd_sc_hd__a32o_1
X_10398_ _10388_/X _10391_/X _10394_/X _10397_/X _11328_/S _11588_/B1 vssd1 vssd1
+ vccd1 vccd1 _10399_/B sky130_fd_sc_hd__mux4_2
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ _12219_/A _12137_/B _12138_/B vssd1 vssd1 vccd1 vccd1 _17840_/D sky130_fd_sc_hd__nor3_1
X_17994_ _19564_/CLK _17994_/D vssd1 vssd1 vccd1 vccd1 _17994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16945_ _18767_/Q _16965_/A2 _16965_/B1 input232/X _16965_/C1 vssd1 vssd1 vccd1 vccd1
+ _16945_/X sky130_fd_sc_hd__a221o_2
X_12068_ _12471_/A0 _12088_/A2 _12067_/X _17328_/A vssd1 vssd1 vccd1 vccd1 _17811_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11019_ _11013_/X _11015_/X _11018_/X _11406_/B2 _09264_/S vssd1 vssd1 vccd1 vccd1
+ _11019_/X sky130_fd_sc_hd__o221a_1
XFILLER_226_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16876_ _16892_/A _16876_/B vssd1 vssd1 vccd1 vccd1 _19303_/D sky130_fd_sc_hd__and2_1
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18615_ _19639_/CLK _18615_/D vssd1 vssd1 vccd1 vccd1 _18615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _18619_/Q _17717_/A0 _15833_/S vssd1 vssd1 vccd1 vccd1 _18619_/D sky130_fd_sc_hd__mux2_1
X_19595_ _19595_/CLK _19595_/D vssd1 vssd1 vccd1 vccd1 _19595_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15758_ _15758_/A _15758_/B vssd1 vssd1 vccd1 vccd1 _15758_/X sky130_fd_sc_hd__xor2_1
X_18546_ _19600_/CLK _18546_/D vssd1 vssd1 vccd1 vccd1 _18546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ _14875_/B1 _14706_/X _14708_/Y _14928_/B1 vssd1 vssd1 vccd1 vccd1 _14710_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_18477_ _19320_/CLK _18477_/D vssd1 vssd1 vccd1 vccd1 _18477_/Q sky130_fd_sc_hd__dfxtp_1
X_15689_ _15689_/A _15689_/B vssd1 vssd1 vccd1 vccd1 _15690_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_390 _17337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17428_ _17428_/A _17462_/B vssd1 vssd1 vccd1 vccd1 _17428_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17359_ _19477_/Q _17184_/B _17361_/S vssd1 vssd1 vccd1 vccd1 _17360_/B sky130_fd_sc_hd__mux2_1
XFILLER_277_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19029_ _19219_/CLK _19029_/D vssd1 vssd1 vccd1 vccd1 _19029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08994_ _08939_/A _08913_/X _08992_/Y vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__a21o_4
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09615_ _09613_/X _09614_/X _10264_/S vssd1 vssd1 vccd1 vccd1 _09615_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09546_ _11172_/A1 _19201_/Q _19169_/Q _09925_/S _11480_/C1 vssd1 vssd1 vccd1 vccd1
+ _09546_/X sky130_fd_sc_hd__a221o_1
XFILLER_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09477_ input167/X input138/X _09990_/S vssd1 vssd1 vccd1 vccd1 _09477_/X sky130_fd_sc_hd__mux2_8
XPHY_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ _12626_/B vssd1 vssd1 vccd1 vccd1 _13387_/A sky130_fd_sc_hd__inv_2
XFILLER_109_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10321_ _10319_/X _10320_/X _11161_/S vssd1 vssd1 vccd1 vccd1 _10321_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ _13354_/A _13039_/X _13038_/Y _13194_/S vssd1 vssd1 vccd1 vccd1 _13040_/X
+ sky130_fd_sc_hd__o211a_1
X_10252_ _18903_/Q _11167_/B _10251_/X _11397_/A1 vssd1 vssd1 vccd1 vccd1 _10252_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10183_ _10334_/A1 _17787_/Q _10090_/S _18336_/Q vssd1 vssd1 vccd1 vccd1 _10183_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_278_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1203 _12754_/Y vssd1 vssd1 vccd1 vccd1 _13962_/B sky130_fd_sc_hd__buf_6
Xfanout1214 _12721_/S vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__buf_6
XFILLER_279_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1225 _15216_/A1 vssd1 vssd1 vccd1 vccd1 _15382_/B2 sky130_fd_sc_hd__buf_4
XFILLER_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14991_ _18500_/Q _15001_/A2 _14990_/Y _14991_/C1 vssd1 vssd1 vccd1 vccd1 _18500_/D
+ sky130_fd_sc_hd__a211o_1
Xfanout1247 _16820_/A3 vssd1 vssd1 vccd1 vccd1 _11216_/A2 sky130_fd_sc_hd__buf_6
Xfanout1258 _13937_/A vssd1 vssd1 vccd1 vccd1 _11441_/B sky130_fd_sc_hd__buf_4
XFILLER_282_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1269 _14591_/A2 vssd1 vssd1 vccd1 vccd1 _14589_/A2 sky130_fd_sc_hd__buf_4
X_16730_ _16737_/A _16730_/B _16736_/D vssd1 vssd1 vccd1 vccd1 _19262_/D sky130_fd_sc_hd__nor3_1
X_13942_ _17854_/Q _13942_/A2 _13942_/B1 _17886_/Q vssd1 vssd1 vccd1 vccd1 _13942_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16661_ _19242_/Q _19241_/Q _16661_/C vssd1 vssd1 vccd1 vccd1 _16667_/C sky130_fd_sc_hd__and3_1
X_13873_ _17948_/Q _13940_/A2 _13872_/X _14029_/C1 vssd1 vssd1 vccd1 vccd1 _17948_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_234_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_175_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19521_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_262_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18400_ _19466_/CLK _18400_/D vssd1 vssd1 vccd1 vccd1 _18400_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15612_ _15612_/A _15612_/B vssd1 vssd1 vccd1 vccd1 _15612_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12824_ _12821_/A _12720_/X _12823_/Y vssd1 vssd1 vccd1 vccd1 _12824_/Y sky130_fd_sc_hd__o21ai_1
X_19380_ _19542_/CLK _19380_/D vssd1 vssd1 vccd1 vccd1 _19380_/Q sky130_fd_sc_hd__dfxtp_1
X_16592_ _16592_/A0 _19195_/Q _16623_/S vssd1 vssd1 vccd1 vccd1 _19195_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_104_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18691_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_222_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18331_ _19638_/CLK _18331_/D vssd1 vssd1 vccd1 vccd1 _18331_/Q sky130_fd_sc_hd__dfxtp_1
X_15543_ _15522_/A _15519_/Y _15521_/B vssd1 vssd1 vccd1 vccd1 _15544_/B sky130_fd_sc_hd__o21a_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12755_ _12755_/A _12756_/B vssd1 vssd1 vccd1 vccd1 _12755_/X sky130_fd_sc_hd__and2_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18262_ _19055_/CLK _18262_/D vssd1 vssd1 vccd1 vccd1 _18262_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11702_/X _11706_/B _11706_/C vssd1 vssd1 vccd1 vccd1 _11706_/X sky130_fd_sc_hd__and3b_4
X_15474_ _15474_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15474_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _09896_/Y _12657_/B _13911_/A vssd1 vssd1 vccd1 vccd1 _12686_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14425_ _18564_/Q _14427_/B vssd1 vssd1 vccd1 vccd1 _18277_/D sky130_fd_sc_hd__and2_1
X_17213_ _17231_/A _17213_/B vssd1 vssd1 vccd1 vccd1 _19422_/D sky130_fd_sc_hd__nor2_1
X_18193_ _19646_/CLK _18193_/D vssd1 vssd1 vccd1 vccd1 _18193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11637_ _11637_/A _13860_/A vssd1 vssd1 vccd1 vccd1 _17531_/A sky130_fd_sc_hd__xor2_4
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17144_ _17255_/A _17144_/B vssd1 vssd1 vccd1 vccd1 _19399_/D sky130_fd_sc_hd__nor2_1
X_14356_ _18208_/Q _17663_/A0 _14380_/S vssd1 vssd1 vccd1 vccd1 _18208_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11568_ _11568_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11568_/X sky130_fd_sc_hd__or2_1
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13307_ _13928_/A1 _13296_/X _13306_/X vssd1 vssd1 vccd1 vccd1 _13998_/B sky130_fd_sc_hd__a21oi_4
X_17075_ _19371_/Q _17113_/B vssd1 vssd1 vccd1 vccd1 _17075_/X sky130_fd_sc_hd__or2_1
X_10519_ _10513_/S _10508_/X _10509_/X vssd1 vssd1 vccd1 vccd1 _10519_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14287_ _11376_/B _18146_/Q _14301_/S vssd1 vssd1 vccd1 vccd1 _18146_/D sky130_fd_sc_hd__mux2_1
X_11499_ _11497_/X _11498_/X _11507_/S vssd1 vssd1 vccd1 vccd1 _11499_/X sky130_fd_sc_hd__mux2_2
XFILLER_109_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16026_ _16020_/Y _16025_/X _16024_/X _16052_/A vssd1 vssd1 vccd1 vccd1 _18727_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13238_ _15303_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13238_/X sky130_fd_sc_hd__and2_1
XFILLER_124_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13169_ _19498_/Q _13064_/B _13243_/B1 _13168_/X vssd1 vssd1 vccd1 vccd1 _13169_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17977_ _18627_/CLK _17977_/D vssd1 vssd1 vccd1 vccd1 _17977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16928_ _16928_/A _16928_/B vssd1 vssd1 vccd1 vccd1 _19316_/D sky130_fd_sc_hd__and2_1
Xfanout1770 _10471_/S vssd1 vssd1 vccd1 vccd1 _11251_/S sky130_fd_sc_hd__buf_6
Xfanout1781 _10373_/S vssd1 vssd1 vccd1 vccd1 _09708_/A sky130_fd_sc_hd__buf_6
XFILLER_284_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1792 _17904_/Q vssd1 vssd1 vccd1 vccd1 _12389_/A1 sky130_fd_sc_hd__buf_12
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19647_ _19647_/CLK _19647_/D vssd1 vssd1 vccd1 vccd1 _19647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16859_ _19299_/Q _16967_/S _16858_/Y _16968_/A vssd1 vssd1 vccd1 vccd1 _19299_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09400_ _09866_/B _15259_/A _09367_/X vssd1 vssd1 vccd1 vccd1 _09401_/C sky130_fd_sc_hd__o21ai_4
XFILLER_53_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19578_ _19638_/CLK _19578_/D vssd1 vssd1 vccd1 vccd1 _19578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09331_ _09331_/A _09331_/B vssd1 vssd1 vccd1 vccd1 _09331_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18529_ _19229_/CLK _18529_/D vssd1 vssd1 vccd1 vccd1 _18529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09262_ _09272_/A1 _19627_/Q _18916_/Q _09252_/S vssd1 vssd1 vccd1 vccd1 _09262_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09193_ _18111_/Q _09367_/B vssd1 vssd1 vccd1 vccd1 _09193_/X sky130_fd_sc_hd__or2_4
XFILLER_119_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08977_ _08977_/A _08977_/B vssd1 vssd1 vccd1 vccd1 _08977_/Y sky130_fd_sc_hd__nor2_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_2_wb_clk_i _19652_/A vssd1 vssd1 vccd1 vccd1 _18613_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10870_ _09107_/D _10859_/X _10867_/X _10869_/X vssd1 vssd1 vccd1 vccd1 _10870_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_244_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09529_ _09527_/X _09528_/X _09935_/A vssd1 vssd1 vccd1 vccd1 _09529_/X sky130_fd_sc_hd__mux2_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ _15857_/A _12506_/X _12534_/X _12539_/X _12510_/X vssd1 vssd1 vccd1 vccd1
+ _12540_/X sky130_fd_sc_hd__o221a_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _12471_/A0 _14675_/B _12482_/S vssd1 vssd1 vccd1 vccd1 _12528_/C sky130_fd_sc_hd__mux2_8
XFILLER_40_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14210_ _14714_/A _14252_/B vssd1 vssd1 vccd1 vccd1 _14210_/Y sky130_fd_sc_hd__nand2_1
X_11422_ _11420_/X _11421_/X _11507_/S vssd1 vssd1 vccd1 vccd1 _11422_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15190_ _19460_/Q _15189_/Y _15400_/S vssd1 vssd1 vccd1 vccd1 _15190_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14141_ _14141_/A _14141_/B _14141_/C _14141_/D vssd1 vssd1 vccd1 vccd1 _14141_/Y
+ sky130_fd_sc_hd__nor4_1
X_11353_ _11594_/A1 _19113_/Q _19145_/Q _11353_/B2 vssd1 vssd1 vccd1 vccd1 _11353_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _11624_/A1 _10239_/B _10303_/X _08957_/Y vssd1 vssd1 vccd1 vccd1 _13843_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14072_ _17722_/A0 _18014_/Q _14072_/S vssd1 vssd1 vccd1 vccd1 _18014_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11284_ _11284_/A1 _18609_/Q _18180_/Q _11284_/B2 vssd1 vssd1 vccd1 vccd1 _11284_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13023_ _13023_/A _13023_/B vssd1 vssd1 vccd1 vccd1 _13023_/X sky130_fd_sc_hd__or2_1
XFILLER_180_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17900_ _18817_/CLK _17900_/D vssd1 vssd1 vccd1 vccd1 _17900_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10235_ _10309_/B _10235_/B vssd1 vssd1 vccd1 vccd1 _10235_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18880_ _18880_/CLK _18880_/D vssd1 vssd1 vccd1 vccd1 _18880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1000 _16618_/A0 vssd1 vssd1 vccd1 vccd1 _17718_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_279_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1011 _15047_/Y vssd1 vssd1 vccd1 vccd1 _15079_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_239_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17831_ _17865_/CLK _17831_/D vssd1 vssd1 vccd1 vccd1 _17831_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1022 _12458_/Y vssd1 vssd1 vccd1 vccd1 _14973_/A1 sky130_fd_sc_hd__buf_4
X_10166_ _17949_/Q _08946_/Y _10165_/X _11451_/B2 vssd1 vssd1 vccd1 vccd1 _10166_/X
+ sky130_fd_sc_hd__o22a_4
Xfanout1033 _16465_/A0 vssd1 vssd1 vccd1 vccd1 _17664_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1044 _08958_/X vssd1 vssd1 vccd1 vccd1 _11055_/B2 sky130_fd_sc_hd__clkbuf_16
Xfanout1055 _15523_/S vssd1 vssd1 vccd1 vccd1 _15781_/S sky130_fd_sc_hd__buf_6
XFILLER_254_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1066 _13486_/A1 vssd1 vssd1 vccd1 vccd1 _13224_/B sky130_fd_sc_hd__buf_2
X_17762_ _19634_/CLK _17762_/D vssd1 vssd1 vccd1 vccd1 _17762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1077 _17659_/A0 vssd1 vssd1 vccd1 vccd1 _16592_/A0 sky130_fd_sc_hd__buf_2
X_10097_ _10243_/A _10096_/Y _10093_/Y _09264_/S vssd1 vssd1 vccd1 vccd1 _10097_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14974_ _14972_/X _14973_/X _14995_/A1 vssd1 vssd1 vccd1 vccd1 _14974_/X sky130_fd_sc_hd__a21o_1
Xfanout1088 _09825_/X vssd1 vssd1 vccd1 vccd1 _16594_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19501_ _19533_/CLK _19501_/D vssd1 vssd1 vccd1 vccd1 _19501_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1099 _08882_/Y vssd1 vssd1 vccd1 vccd1 _17516_/C1 sky130_fd_sc_hd__buf_4
XFILLER_235_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16713_ _19257_/Q _19256_/Q _16713_/C vssd1 vssd1 vccd1 vccd1 _16715_/B sky130_fd_sc_hd__and3_1
XFILLER_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ _19390_/Q _13924_/X _13925_/S vssd1 vssd1 vccd1 vccd1 _13925_/X sky130_fd_sc_hd__mux2_1
XFILLER_267_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17693_ _17693_/A0 _19619_/Q _17719_/S vssd1 vssd1 vccd1 vccd1 _19619_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19432_ _19433_/CLK _19432_/D vssd1 vssd1 vccd1 vccd1 _19432_/Q sky130_fd_sc_hd__dfxtp_1
X_16644_ _16740_/A _16649_/C vssd1 vssd1 vccd1 vccd1 _16644_/Y sky130_fd_sc_hd__nor2_1
X_13856_ _14030_/B vssd1 vssd1 vccd1 vccd1 _13856_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12807_ _12803_/Y _12806_/X _13130_/A vssd1 vssd1 vccd1 vccd1 _12807_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19363_ _19363_/CLK _19363_/D vssd1 vssd1 vccd1 vccd1 _19363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13787_ _13928_/A1 _13776_/X _13778_/Y _13786_/Y vssd1 vssd1 vccd1 vccd1 _14026_/B
+ sky130_fd_sc_hd__o2bb2a_4
X_16575_ _16608_/A0 _19179_/Q _16586_/S vssd1 vssd1 vccd1 vccd1 _19179_/D sky130_fd_sc_hd__mux2_1
X_10999_ _18034_/Q _18002_/Q _11386_/S vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18314_ _19614_/CLK _18314_/D vssd1 vssd1 vccd1 vccd1 _18314_/Q sky130_fd_sc_hd__dfxtp_1
X_12738_ _13414_/A _12737_/X _12719_/X vssd1 vssd1 vccd1 vccd1 _12738_/Y sky130_fd_sc_hd__o21ai_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15526_ _15526_/A _15526_/B vssd1 vssd1 vccd1 vccd1 _15526_/Y sky130_fd_sc_hd__nor2_1
X_19294_ _19327_/CLK _19294_/D vssd1 vssd1 vccd1 vccd1 _19294_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18245_ _19627_/CLK _18245_/D vssd1 vssd1 vccd1 vccd1 _18245_/Q sky130_fd_sc_hd__dfxtp_1
X_15457_ _15457_/A vssd1 vssd1 vccd1 vccd1 _15457_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12669_ _09143_/A _10908_/B _13911_/A vssd1 vssd1 vccd1 vccd1 _12669_/X sky130_fd_sc_hd__mux2_2
XFILLER_204_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14408_ _17715_/A0 _18259_/Q _14416_/S vssd1 vssd1 vccd1 vccd1 _18259_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18176_ _19629_/CLK _18176_/D vssd1 vssd1 vccd1 vccd1 _18176_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_72_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18543_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15388_ _18575_/Q _18574_/Q _15388_/C vssd1 vssd1 vccd1 vccd1 _15412_/B sky130_fd_sc_hd__and3_1
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14339_ _18196_/Q _16292_/A0 _14339_/S vssd1 vssd1 vccd1 vccd1 _18196_/D sky130_fd_sc_hd__mux2_1
X_17127_ _15118_/Y _17120_/Y _17404_/A _17141_/A vssd1 vssd1 vccd1 vccd1 _17127_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_274_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ _17563_/A _17114_/A2 _17057_/X _17378_/A vssd1 vssd1 vccd1 vccd1 _19362_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16009_ _18720_/Q _16019_/A2 _16008_/X _16153_/D vssd1 vssd1 vccd1 vccd1 _18720_/D
+ sky130_fd_sc_hd__o211a_1
X_08900_ _10663_/S _12442_/B vssd1 vssd1 vccd1 vccd1 _08900_/Y sky130_fd_sc_hd__nand2_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09878_/X _09879_/X _11189_/A vssd1 vssd1 vccd1 vccd1 _09880_/X sky130_fd_sc_hd__mux2_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _18132_/Q vssd1 vssd1 vccd1 vccd1 _14268_/A sky130_fd_sc_hd__clkinv_4
XFILLER_253_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09314_ _09946_/B1 _15284_/A _09281_/Y vssd1 vssd1 vccd1 vccd1 _09317_/B sky130_fd_sc_hd__o21ai_4
XFILLER_179_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09245_ _09245_/A _11556_/B _09245_/C _09245_/D vssd1 vssd1 vccd1 vccd1 _09903_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09176_ _09174_/X _09175_/X _09264_/S vssd1 vssd1 vccd1 vccd1 _09176_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10020_ _11251_/S _10020_/B _10020_/C vssd1 vssd1 vccd1 vccd1 _10020_/X sky130_fd_sc_hd__and3_1
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput103 dout0[6] vssd1 vssd1 vccd1 vccd1 input103/X sky130_fd_sc_hd__clkbuf_2
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput114 dout1[16] vssd1 vssd1 vccd1 vccd1 input114/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput125 dout1[26] vssd1 vssd1 vccd1 vccd1 input125/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 dout1[36] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_hd__buf_2
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput147 dout1[46] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput158 dout1[56] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_hd__buf_2
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput169 dout1[8] vssd1 vssd1 vccd1 vccd1 input169/X sky130_fd_sc_hd__clkbuf_2
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _18734_/Q _18733_/Q vssd1 vssd1 vccd1 vccd1 _11972_/D sky130_fd_sc_hd__nand2_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _17943_/Q _13742_/A2 _13709_/X _14417_/A vssd1 vssd1 vccd1 vccd1 _17943_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10922_ _18426_/Q _11300_/B _10921_/X _10784_/S vssd1 vssd1 vccd1 vccd1 _10922_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_260_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _16819_/B _15834_/B vssd1 vssd1 vccd1 vccd1 _14690_/Y sky130_fd_sc_hd__nor2_4
XFILLER_17_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13641_ _18122_/Q _13642_/B vssd1 vssd1 vccd1 vccd1 _13704_/C sky130_fd_sc_hd__and2_2
X_10853_ _19638_/Q _18927_/Q _10853_/S vssd1 vssd1 vccd1 vccd1 _10853_/X sky130_fd_sc_hd__mux2_1
XFILLER_260_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16592_/A0 _18971_/Q _16391_/S vssd1 vssd1 vccd1 vccd1 _18971_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13572_ _13602_/B2 _13313_/X _13315_/X _12704_/S vssd1 vssd1 vccd1 vccd1 _13572_/X
+ sky130_fd_sc_hd__o22a_1
X_10784_ _10782_/X _10783_/X _10784_/S vssd1 vssd1 vccd1 vccd1 _10785_/B sky130_fd_sc_hd__mux2_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _15365_/C _15312_/B vssd1 vssd1 vccd1 vccd1 _15313_/A sky130_fd_sc_hd__or2_1
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12523_ _12577_/A _12578_/A vssd1 vssd1 vccd1 vccd1 _12768_/B sky130_fd_sc_hd__or2_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _16622_/A0 _18905_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _18905_/D sky130_fd_sc_hd__mux2_1
XFILLER_169_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18030_ _18613_/CLK _18030_/D vssd1 vssd1 vccd1 vccd1 _18030_/Q sky130_fd_sc_hd__dfxtp_1
X_15242_ _14220_/A _15786_/A2 _15239_/Y _12318_/A _15243_/B vssd1 vssd1 vccd1 vccd1
+ _15242_/X sky130_fd_sc_hd__o221a_1
X_12454_ _12455_/A _12587_/B vssd1 vssd1 vccd1 vccd1 _12454_/X sky130_fd_sc_hd__and2_2
XFILLER_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11405_ _11403_/X _11404_/X _11481_/A vssd1 vssd1 vccd1 vccd1 _11405_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15173_ _15173_/A _15259_/B vssd1 vssd1 vccd1 vccd1 _15173_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ _17887_/Q _12433_/B _12385_/C vssd1 vssd1 vccd1 vccd1 _12385_/X sky130_fd_sc_hd__or3_1
XFILLER_67_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14124_ _17674_/A0 _18063_/Q _14131_/S vssd1 vssd1 vccd1 vccd1 _18063_/D sky130_fd_sc_hd__mux2_1
X_11336_ _12596_/A vssd1 vssd1 vccd1 vccd1 _11368_/A sky130_fd_sc_hd__inv_2
XFILLER_126_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14055_ _17672_/A0 _17997_/Q _14070_/S vssd1 vssd1 vccd1 vccd1 _17997_/D sky130_fd_sc_hd__mux2_1
X_18932_ _19643_/CLK _18932_/D vssd1 vssd1 vccd1 vccd1 _18932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11267_ _11282_/A _11262_/X _11266_/X vssd1 vssd1 vccd1 vccd1 _11267_/Y sky130_fd_sc_hd__a21oi_1
X_13006_ _17924_/Q _13808_/C1 _13005_/X vssd1 vssd1 vccd1 vccd1 _13007_/B sky130_fd_sc_hd__a21oi_1
XFILLER_279_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10218_ _18872_/Q _10215_/S _10293_/B1 vssd1 vssd1 vccd1 vccd1 _10218_/X sky130_fd_sc_hd__o21a_1
X_18863_ _19055_/CLK _18863_/D vssd1 vssd1 vccd1 vccd1 _18863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11198_ _11196_/X _11197_/X _11198_/S vssd1 vssd1 vccd1 vccd1 _11198_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_190_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19609_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17814_ _17814_/CLK _17814_/D vssd1 vssd1 vccd1 vccd1 _17814_/Q sky130_fd_sc_hd__dfxtp_4
X_10149_ _18469_/Q _18370_/Q _10206_/S vssd1 vssd1 vccd1 vccd1 _10149_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18794_ _19025_/CLK _18794_/D vssd1 vssd1 vccd1 vccd1 _18794_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17745_ _18645_/Q vssd1 vssd1 vccd1 vccd1 _18645_/D sky130_fd_sc_hd__clkbuf_2
X_14957_ input61/X input96/X _15007_/S vssd1 vssd1 vccd1 vccd1 _14958_/A sky130_fd_sc_hd__mux2_2
XFILLER_94_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _13908_/A _13908_/B vssd1 vssd1 vccd1 vccd1 _14152_/C sky130_fd_sc_hd__xnor2_4
XFILLER_251_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17676_ _17676_/A0 _19603_/Q _17690_/S vssd1 vssd1 vccd1 vccd1 _19603_/D sky130_fd_sc_hd__mux2_1
X_14888_ _14979_/A1 _18271_/Q _14887_/Y _14918_/B1 vssd1 vssd1 vccd1 vccd1 _14888_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_90_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19415_ _19482_/CLK _19415_/D vssd1 vssd1 vccd1 vccd1 _19415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16627_ _19230_/Q input250/X _16627_/S vssd1 vssd1 vccd1 vccd1 _19230_/D sky130_fd_sc_hd__mux2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13839_ _13899_/A _13835_/X _13838_/X _13869_/B2 vssd1 vssd1 vccd1 vccd1 _13839_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_251_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19346_ _19540_/CLK _19346_/D vssd1 vssd1 vccd1 vccd1 _19346_/Q sky130_fd_sc_hd__dfxtp_1
X_16558_ _17625_/A _16591_/B vssd1 vssd1 vccd1 vccd1 _16558_/Y sky130_fd_sc_hd__nand2_2
XFILLER_188_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15509_ _15508_/B _15489_/B _15482_/Y vssd1 vssd1 vccd1 vccd1 _15511_/B sky130_fd_sc_hd__a21oi_1
X_19277_ _19280_/CLK _19277_/D vssd1 vssd1 vccd1 vccd1 _19277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16489_ _16522_/A0 _19096_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _19096_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09030_ _09025_/A _09025_/B _09986_/B _10085_/A vssd1 vssd1 vccd1 vccd1 _09030_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_176_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18228_ _19649_/CLK _18228_/D vssd1 vssd1 vccd1 vccd1 _18228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18159_ _19055_/CLK _18159_/D vssd1 vssd1 vccd1 vccd1 _18159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09932_ _19196_/Q _19164_/Q _11472_/C vssd1 vssd1 vccd1 vccd1 _09932_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout804 _16161_/Y vssd1 vssd1 vccd1 vccd1 _16165_/S sky130_fd_sc_hd__buf_12
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout815 _14380_/S vssd1 vssd1 vccd1 vccd1 _14382_/S sky130_fd_sc_hd__buf_12
XFILLER_258_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout826 _11990_/Y vssd1 vssd1 vccd1 vccd1 _12022_/S sky130_fd_sc_hd__buf_12
XFILLER_98_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09863_ _12320_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _09863_/Y sky130_fd_sc_hd__nand2_2
Xfanout837 _11067_/X vssd1 vssd1 vccd1 vccd1 _16543_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout848 _14510_/A0 vssd1 vssd1 vccd1 vccd1 _17679_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_259_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout859 _10682_/X vssd1 vssd1 vccd1 vccd1 _10713_/A2 sky130_fd_sc_hd__buf_4
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09792_/X _09793_/X _10040_/S vssd1 vssd1 vccd1 vccd1 _09794_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _18564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_219 _18626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09228_ _12599_/A _09229_/B vssd1 vssd1 vccd1 vccd1 _13230_/S sky130_fd_sc_hd__nor2_1
XFILLER_155_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09159_ _11687_/A _09157_/X _09158_/X vssd1 vssd1 vccd1 vccd1 _09159_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12170_ _17853_/Q _12170_/B vssd1 vssd1 vccd1 vccd1 _12176_/C sky130_fd_sc_hd__and2_2
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11121_ _18860_/Q _18892_/Q _19052_/Q _19020_/Q _11125_/B2 _11338_/S1 vssd1 vssd1
+ vccd1 vccd1 _11121_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11052_ _11028_/Y _11032_/Y _11438_/B1 vssd1 vssd1 vccd1 vccd1 _11052_/X sky130_fd_sc_hd__a21o_1
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10003_ _11567_/S _10001_/X _10002_/X _09853_/S vssd1 vssd1 vccd1 vccd1 _10003_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_277_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15860_ _15860_/A _15905_/B _15908_/C vssd1 vssd1 vccd1 vccd1 _15860_/X sky130_fd_sc_hd__and3_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14811_ _18113_/Q _14994_/B vssd1 vssd1 vccd1 vccd1 _14811_/X sky130_fd_sc_hd__or2_1
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _18593_/Q _15791_/B vssd1 vssd1 vccd1 vccd1 _15791_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _19517_/Q _17517_/B _17529_/X vssd1 vssd1 vccd1 vccd1 _19517_/D sky130_fd_sc_hd__o21ba_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _14992_/A1 _13024_/X _14973_/B1 _18631_/Q _14741_/B vssd1 vssd1 vccd1 vccd1
+ _14742_/X sky130_fd_sc_hd__a221o_1
XFILLER_18_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11954_ _11666_/A _11774_/X _11663_/A vssd1 vssd1 vccd1 vccd1 _14343_/C sky130_fd_sc_hd__a21o_1
XFILLER_91_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _18121_/Q _10904_/Y _10905_/S vssd1 vssd1 vccd1 vccd1 _10908_/B sky130_fd_sc_hd__mux2_4
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14673_ _14688_/B _14680_/B _14680_/C _14672_/C vssd1 vssd1 vccd1 vccd1 _14673_/X
+ sky130_fd_sc_hd__or4b_1
X_17461_ _18576_/Q _17461_/A2 _17460_/X _17546_/A2 vssd1 vssd1 vccd1 vccd1 _17461_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_199_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11885_ _11811_/Y _11875_/Y _11884_/X vssd1 vssd1 vccd1 vccd1 _11886_/C sky130_fd_sc_hd__o21ai_2
XFILLER_233_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19200_ _19653_/A _19200_/D vssd1 vssd1 vccd1 vccd1 _19200_/Q sky130_fd_sc_hd__dfxtp_1
X_16412_ _16610_/A0 _19021_/Q _16424_/S vssd1 vssd1 vccd1 vccd1 _19021_/D sky130_fd_sc_hd__mux2_1
X_13624_ _17844_/Q _13744_/A2 _13744_/B1 _17876_/Q vssd1 vssd1 vccd1 vccd1 _13624_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10836_ _11143_/A1 _10834_/Y _10835_/X vssd1 vssd1 vccd1 vccd1 _10836_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17392_ _14424_/A _17391_/X _17437_/A2 _18777_/Q vssd1 vssd1 vccd1 vccd1 _17392_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_198_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19131_ _19195_/CLK _19131_/D vssd1 vssd1 vccd1 vccd1 _19131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16343_ _18955_/Q _16542_/A0 _16352_/S vssd1 vssd1 vccd1 vccd1 _18955_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13555_ _19411_/Q _13948_/A2 _13948_/B1 vssd1 vssd1 vccd1 vccd1 _13555_/X sky130_fd_sc_hd__a21o_1
XFILLER_160_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10767_ _10763_/X _10766_/X _11328_/S vssd1 vssd1 vccd1 vccd1 _10767_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12506_ _13167_/A _13165_/B vssd1 vssd1 vccd1 vccd1 _12506_/X sky130_fd_sc_hd__or2_4
XFILLER_160_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16274_ _11376_/B _18888_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _18888_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19062_ _19645_/CLK _19062_/D vssd1 vssd1 vccd1 vccd1 _19062_/Q sky130_fd_sc_hd__dfxtp_1
X_13486_ _13486_/A1 _14146_/B _13909_/B1 vssd1 vssd1 vccd1 vccd1 _13486_/Y sky130_fd_sc_hd__a21oi_1
X_10698_ _18554_/Q _18429_/Q _18038_/Q _18006_/Q _11249_/S _11156_/C1 vssd1 vssd1
+ vccd1 vccd1 _10698_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18013_ _19615_/CLK _18013_/D vssd1 vssd1 vccd1 vccd1 _18013_/Q sky130_fd_sc_hd__dfxtp_1
X_15225_ _18567_/Q _15224_/C _18568_/Q vssd1 vssd1 vccd1 vccd1 _15226_/B sky130_fd_sc_hd__a21oi_1
X_12437_ _12437_/A _12587_/B vssd1 vssd1 vccd1 vccd1 _12437_/Y sky130_fd_sc_hd__nand2_1
Xoutput407 _11929_/X vssd1 vssd1 vccd1 vccd1 din0[9] sky130_fd_sc_hd__buf_4
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15156_ _15171_/A _15156_/B vssd1 vssd1 vccd1 vccd1 _15156_/X sky130_fd_sc_hd__and2_1
Xoutput418 _18488_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[17] sky130_fd_sc_hd__buf_4
X_12368_ _17897_/Q _12408_/B _12367_/Y _13981_/C1 vssd1 vssd1 vccd1 vccd1 _17897_/D
+ sky130_fd_sc_hd__o211a_1
Xoutput429 _18498_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[27] sky130_fd_sc_hd__buf_4
XFILLER_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14107_ _17690_/A0 _18047_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _18047_/D sky130_fd_sc_hd__mux2_1
XFILLER_259_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11319_ _11327_/S _11572_/A1 _19209_/Q _11578_/S vssd1 vssd1 vccd1 vccd1 _11319_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15087_ _19390_/Q _15088_/B _15087_/C vssd1 vssd1 vccd1 vccd1 _15101_/A sky130_fd_sc_hd__and3_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12299_ _18082_/Q _18081_/Q _12277_/B vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__or3b_4
XFILLER_113_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18915_ _19626_/CLK _18915_/D vssd1 vssd1 vccd1 vccd1 _18915_/Q sky130_fd_sc_hd__dfxtp_1
X_14038_ _17800_/Q _16392_/B _16392_/C vssd1 vssd1 vccd1 vccd1 _17658_/A sky130_fd_sc_hd__and3b_4
XFILLER_268_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18846_ _19589_/CLK _18846_/D vssd1 vssd1 vccd1 vccd1 _18846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18777_ _18778_/CLK _18777_/D vssd1 vssd1 vccd1 vccd1 _18777_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_283_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15989_ _18710_/Q _16005_/A2 _15988_/X _14203_/A vssd1 vssd1 vccd1 vccd1 _18710_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17728_ _18628_/Q vssd1 vssd1 vccd1 vccd1 _18628_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17659_ _17659_/A0 _19586_/Q _17681_/S vssd1 vssd1 vccd1 vccd1 _19586_/D sky130_fd_sc_hd__mux2_1
XFILLER_224_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19329_ _19522_/CLK _19329_/D vssd1 vssd1 vccd1 vccd1 _19329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ _09245_/A _09031_/S vssd1 vssd1 vccd1 vccd1 _09013_/Y sky130_fd_sc_hd__nor2_2
XFILLER_275_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout601 _17724_/B vssd1 vssd1 vccd1 vccd1 _14244_/B sky130_fd_sc_hd__buf_8
Xfanout612 _11799_/A vssd1 vssd1 vccd1 vccd1 _11926_/A1 sky130_fd_sc_hd__buf_8
XFILLER_259_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09915_ _11404_/A1 _17759_/Q _11481_/C _18308_/Q _09935_/A vssd1 vssd1 vccd1 vccd1
+ _09915_/X sky130_fd_sc_hd__o221a_1
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout623 _16980_/X vssd1 vssd1 vccd1 vccd1 _17032_/A2 sky130_fd_sc_hd__buf_6
XFILLER_101_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout634 _11826_/A vssd1 vssd1 vccd1 vccd1 _11859_/B sky130_fd_sc_hd__buf_8
Xfanout645 _17050_/X vssd1 vssd1 vccd1 vccd1 _17074_/A2 sky130_fd_sc_hd__buf_4
Xfanout656 _13277_/S vssd1 vssd1 vccd1 vccd1 _13372_/S sky130_fd_sc_hd__buf_6
XFILLER_259_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout667 _11859_/A vssd1 vssd1 vccd1 vccd1 _11820_/A sky130_fd_sc_hd__clkbuf_16
X_09846_ _09854_/A _18206_/Q _12023_/A vssd1 vssd1 vccd1 vccd1 _09846_/X sky130_fd_sc_hd__or3_1
Xfanout678 _12566_/Y vssd1 vssd1 vccd1 vccd1 _13246_/B1 sky130_fd_sc_hd__buf_6
XFILLER_100_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout689 _13244_/B1 vssd1 vssd1 vccd1 vccd1 _13654_/B1 sky130_fd_sc_hd__buf_4
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09777_ _09777_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _09777_/Y sky130_fd_sc_hd__nand2_2
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11670_ _13676_/B vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__clkinv_2
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10621_ _10619_/X _10620_/X _10866_/S vssd1 vssd1 vccd1 vccd1 _10621_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13340_ _19373_/Q _13339_/X _13925_/S vssd1 vssd1 vccd1 vccd1 _13340_/X sky130_fd_sc_hd__mux2_2
XFILLER_139_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ _10550_/X _10551_/X _10784_/S vssd1 vssd1 vccd1 vccd1 _10552_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13271_ _18112_/Q _18111_/Q _13271_/C vssd1 vssd1 vccd1 vccd1 _13326_/B sky130_fd_sc_hd__and3_1
XFILLER_155_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10483_ _10707_/A _10483_/B vssd1 vssd1 vccd1 vccd1 _10483_/X sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_129_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19464_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15010_ _15006_/Y _15009_/X _15010_/B1 vssd1 vssd1 vccd1 vccd1 _15010_/Y sky130_fd_sc_hd__a21oi_4
X_12222_ _17872_/Q _12224_/C _12221_/Y vssd1 vssd1 vccd1 vccd1 _17872_/D sky130_fd_sc_hd__o21a_1
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12153_ _17159_/A _12153_/B _12154_/B vssd1 vssd1 vccd1 vccd1 _17846_/D sky130_fd_sc_hd__nor3_1
XFILLER_162_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11104_ _08874_/D _11135_/S _11181_/B1 _11103_/Y vssd1 vssd1 vccd1 vccd1 _11138_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16961_ _18771_/Q _16961_/A2 _16969_/B1 input236/X _16969_/C1 vssd1 vssd1 vccd1 vccd1
+ _16961_/X sky130_fd_sc_hd__a221o_1
X_12084_ _17917_/Q _12088_/A2 _12083_/X _17328_/A vssd1 vssd1 vccd1 vccd1 _17819_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18700_ _18700_/CLK _18700_/D vssd1 vssd1 vccd1 vccd1 _18700_/Q sky130_fd_sc_hd__dfxtp_1
X_11035_ _11506_/A1 _18957_/Q _18222_/Q _11426_/B2 vssd1 vssd1 vccd1 vccd1 _11035_/X
+ sky130_fd_sc_hd__a22o_1
X_15912_ _18679_/Q _15918_/A2 _15945_/C1 _15911_/X vssd1 vssd1 vccd1 vccd1 _15912_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_238_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16892_ _16892_/A _16892_/B vssd1 vssd1 vccd1 vccd1 _19307_/D sky130_fd_sc_hd__and2_1
XFILLER_231_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18631_ _19622_/CLK _18631_/D vssd1 vssd1 vccd1 vccd1 _18631_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _15843_/A _15843_/B vssd1 vssd1 vccd1 vccd1 _15843_/Y sky130_fd_sc_hd__nand2_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18562_ _19126_/CLK _18562_/D vssd1 vssd1 vccd1 vccd1 _18562_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _15623_/A _15770_/Y _15773_/X vssd1 vssd1 vccd1 vccd1 _15774_/X sky130_fd_sc_hd__a21o_1
X_12986_ _11737_/X _13312_/A _13260_/A vssd1 vssd1 vccd1 vccd1 _12986_/X sky130_fd_sc_hd__o21a_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _17513_/A _17523_/B vssd1 vssd1 vccd1 vccd1 _17513_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _14913_/B1 _14723_/X _14724_/X _14690_/Y vssd1 vssd1 vccd1 vccd1 _14725_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18493_ _19286_/CLK _18493_/D vssd1 vssd1 vccd1 vccd1 _18493_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11937_ _11959_/B2 _11844_/B _11945_/B1 input223/X vssd1 vssd1 vccd1 vccd1 _11937_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _19500_/Q _17453_/B _17442_/X _17443_/Y _17338_/A vssd1 vssd1 vccd1 vccd1
+ _19500_/D sky130_fd_sc_hd__o221a_1
X_14656_ _16615_/A0 _18462_/Q _14664_/S vssd1 vssd1 vccd1 vccd1 _18462_/D sky130_fd_sc_hd__mux2_1
X_11868_ _11909_/A _11868_/B vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__and2_1
XFILLER_159_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10819_ _11601_/A _10814_/X _10818_/X _11602_/C1 vssd1 vssd1 vccd1 vccd1 _10819_/X
+ sky130_fd_sc_hd__o211a_1
X_13607_ _18120_/Q _13606_/C _18121_/Q vssd1 vssd1 vccd1 vccd1 _13608_/B sky130_fd_sc_hd__a21oi_1
XFILLER_220_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17375_ _19485_/Q _17208_/B _17379_/S vssd1 vssd1 vccd1 vccd1 _17376_/B sky130_fd_sc_hd__mux2_1
XFILLER_158_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14587_ _18402_/Q _14589_/A2 _14589_/B1 input31/X vssd1 vssd1 vccd1 vccd1 _14588_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11799_ _11799_/A _11799_/B _11865_/B vssd1 vssd1 vccd1 vccd1 _11799_/X sky130_fd_sc_hd__and3_1
X_19114_ _19114_/CLK _19114_/D vssd1 vssd1 vccd1 vccd1 _19114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16326_ _16326_/A _16459_/C vssd1 vssd1 vccd1 vccd1 _16326_/Y sky130_fd_sc_hd__nor2_8
X_13538_ _13531_/Y _13534_/Y _13537_/X _13966_/C1 vssd1 vssd1 vccd1 vccd1 _13538_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19045_ _19594_/CLK _19045_/D vssd1 vssd1 vccd1 vccd1 _19045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16257_ _16621_/A0 _18872_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _18872_/D sky130_fd_sc_hd__mux2_1
X_13469_ _13962_/B _13468_/X _11215_/B vssd1 vssd1 vccd1 vccd1 _13469_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15208_ _12788_/B _15207_/Y _15307_/B vssd1 vssd1 vccd1 vccd1 _15208_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16188_ _17718_/A0 _18805_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _18805_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ _18564_/Q _15369_/A _15138_/X _15140_/B vssd1 vssd1 vccd1 vccd1 _15139_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _18847_/Q _18879_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09700_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09631_ _10323_/A1 _19200_/Q _19168_/Q _10313_/S _11480_/C1 vssd1 vssd1 vccd1 vccd1
+ _09631_/X sky130_fd_sc_hd__a221o_1
XFILLER_283_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18829_ _19075_/CLK _18829_/D vssd1 vssd1 vccd1 vccd1 _18829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09562_ _18106_/Q _09948_/B vssd1 vssd1 vccd1 vccd1 _09562_/X sky130_fd_sc_hd__or2_1
XFILLER_237_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09493_ _11190_/A1 _19201_/Q _19169_/Q _09952_/S _12766_/A0 vssd1 vssd1 vccd1 vccd1
+ _09493_/X sky130_fd_sc_hd__a221o_1
XFILLER_270_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1407 _09092_/Y vssd1 vssd1 vccd1 vccd1 fanout1407/X sky130_fd_sc_hd__buf_4
Xfanout1418 _09252_/S vssd1 vssd1 vccd1 vccd1 _09269_/S sky130_fd_sc_hd__buf_6
XFILLER_48_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1429 _10326_/A vssd1 vssd1 vccd1 vccd1 _10399_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_171_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout497 _11949_/B1 vssd1 vssd1 vccd1 vccd1 _11945_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09829_ _09853_/S _09829_/B vssd1 vssd1 vccd1 vccd1 _09829_/X sky130_fd_sc_hd__and2_1
XFILLER_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _12440_/X _13911_/B _12835_/Y _12839_/X _14153_/A vssd1 vssd1 vccd1 vccd1
+ _12840_/X sky130_fd_sc_hd__a2111o_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12771_/A _13277_/S vssd1 vssd1 vccd1 vccd1 _12771_/X sky130_fd_sc_hd__or2_4
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11718_/Y _11719_/X _11721_/Y vssd1 vssd1 vccd1 vccd1 _11722_/X sky130_fd_sc_hd__a21o_1
X_14510_ _14510_/A0 _18360_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _18360_/D sky130_fd_sc_hd__mux2_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15789_/A1 _15489_/Y _15537_/B1 vssd1 vssd1 vccd1 vccd1 _15490_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _18580_/Q _14452_/B vssd1 vssd1 vccd1 vccd1 _18293_/D sky130_fd_sc_hd__and2_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11653_ _11653_/A _11653_/B vssd1 vssd1 vccd1 vccd1 _11818_/A sky130_fd_sc_hd__or2_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10604_ _13727_/A vssd1 vssd1 vccd1 vccd1 _10604_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14372_ _18224_/Q _17679_/A0 _14383_/S vssd1 vssd1 vccd1 vccd1 _18224_/D sky130_fd_sc_hd__mux2_1
X_17160_ _17166_/A _17585_/A vssd1 vssd1 vccd1 vccd1 _17457_/A sky130_fd_sc_hd__nand2_1
XFILLER_155_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11584_ _11584_/A1 _19649_/Q _18938_/Q _11302_/S _11584_/C1 vssd1 vssd1 vccd1 vccd1
+ _11584_/X sky130_fd_sc_hd__a221o_1
XFILLER_156_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16111_ _18758_/Q _16137_/B vssd1 vssd1 vccd1 vccd1 _16111_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13323_ _15426_/B _13323_/B vssd1 vssd1 vccd1 vccd1 _13323_/X sky130_fd_sc_hd__or2_4
XFILLER_182_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10535_ _10533_/X _10534_/X _10618_/S vssd1 vssd1 vccd1 vccd1 _10536_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17091_ _19379_/Q _17115_/B vssd1 vssd1 vccd1 vccd1 _17091_/X sky130_fd_sc_hd__or2_1
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16042_ _16039_/X _16041_/X _15845_/A vssd1 vssd1 vccd1 vccd1 _16051_/S sky130_fd_sc_hd__a21o_4
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13254_ _13462_/A _13252_/X _13253_/Y _13224_/A _13254_/B2 vssd1 vssd1 vccd1 vccd1
+ _13255_/B sky130_fd_sc_hd__a32o_1
XFILLER_171_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ _18261_/Q _18836_/Q _10467_/S vssd1 vssd1 vccd1 vccd1 _10466_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12205_ _17866_/Q _12208_/C _16811_/A vssd1 vssd1 vccd1 vccd1 _12205_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _13185_/A _13185_/B _13185_/C _13185_/D vssd1 vssd1 vccd1 vccd1 _13185_/X
+ sky130_fd_sc_hd__or4_1
X_10397_ _10395_/X _10396_/X _10866_/S vssd1 vssd1 vccd1 vccd1 _10397_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12136_ _17839_/Q _17840_/Q _12136_/C vssd1 vssd1 vccd1 vccd1 _12138_/B sky130_fd_sc_hd__and3_1
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17993_ _19595_/CLK _17993_/D vssd1 vssd1 vccd1 vccd1 _17993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16944_ _16960_/A _16944_/B vssd1 vssd1 vccd1 vccd1 _19320_/D sky130_fd_sc_hd__and2_1
XFILLER_150_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12067_ _17811_/Q _12087_/B vssd1 vssd1 vccd1 vccd1 _12067_/X sky130_fd_sc_hd__or2_1
XFILLER_78_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_97_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19076_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11018_ _11016_/X _11017_/X _11481_/A vssd1 vssd1 vccd1 vccd1 _11018_/X sky130_fd_sc_hd__mux2_1
X_16875_ _19303_/Q _17573_/A _16971_/S vssd1 vssd1 vccd1 vccd1 _16876_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19133_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18614_ _19219_/CLK _18614_/D vssd1 vssd1 vccd1 vccd1 _18614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _18618_/Q _17716_/A0 _15833_/S vssd1 vssd1 vccd1 vccd1 _18618_/D sky130_fd_sc_hd__mux2_1
X_19594_ _19594_/CLK _19594_/D vssd1 vssd1 vccd1 vccd1 _19594_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18545_ _19599_/CLK _18545_/D vssd1 vssd1 vccd1 vccd1 _18545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _15757_/A _15757_/B vssd1 vssd1 vccd1 vccd1 _15758_/B sky130_fd_sc_hd__nand2_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _19494_/Q _13064_/B _13243_/B1 _12968_/X vssd1 vssd1 vccd1 vccd1 _12969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_240_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14708_ _14718_/A _14708_/B vssd1 vssd1 vccd1 vccd1 _14708_/Y sky130_fd_sc_hd__nor2_1
X_18476_ _19320_/CLK _18476_/D vssd1 vssd1 vccd1 vccd1 _18476_/Q sky130_fd_sc_hd__dfxtp_1
X_15688_ _15644_/B _15686_/X _15725_/B _15744_/A vssd1 vssd1 vccd1 vccd1 _15689_/B
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_380 _14978_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_391 _08887_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17427_ _18108_/Q _17437_/A2 _17425_/X _17426_/X vssd1 vssd1 vccd1 vccd1 _17427_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14639_ _17665_/A0 _18445_/Q _14660_/S vssd1 vssd1 vccd1 vccd1 _18445_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17358_ _17376_/A _17358_/B vssd1 vssd1 vccd1 vccd1 _19476_/D sky130_fd_sc_hd__and2_1
XFILLER_119_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16309_ _17707_/A0 _18922_/Q _16320_/S vssd1 vssd1 vccd1 vccd1 _18922_/D sky130_fd_sc_hd__mux2_1
X_17289_ _19447_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17289_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19028_ _19609_/CLK _19028_/D vssd1 vssd1 vccd1 vccd1 _19028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08993_ _08939_/A _08913_/X _08992_/Y vssd1 vssd1 vccd1 vccd1 _11556_/B sky130_fd_sc_hd__a21oi_4
XFILLER_130_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09614_ _10323_/A1 _17763_/Q _10313_/S _18312_/Q vssd1 vssd1 vccd1 vccd1 _09614_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09545_ _19041_/Q _19009_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _09545_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09476_ _18107_/Q _09948_/B vssd1 vssd1 vccd1 vccd1 _09476_/X sky130_fd_sc_hd__or2_1
XPHY_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _18621_/Q _18192_/Q _10320_/S vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10251_ _18871_/Q _10253_/C vssd1 vssd1 vccd1 vccd1 _10251_/X sky130_fd_sc_hd__or2_1
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10182_ _10334_/A1 _19583_/Q _10090_/S _19615_/Q vssd1 vssd1 vccd1 vccd1 _10182_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_182_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1204 _12754_/Y vssd1 vssd1 vccd1 vccd1 _13358_/A1 sky130_fd_sc_hd__buf_4
XFILLER_278_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1215 _13863_/B2 vssd1 vssd1 vccd1 vccd1 _13896_/B2 sky130_fd_sc_hd__buf_6
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1226 _12314_/X vssd1 vssd1 vccd1 vccd1 _15216_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1237 _09899_/X vssd1 vssd1 vccd1 vccd1 _11371_/B1 sky130_fd_sc_hd__buf_4
X_14990_ _14986_/Y _14989_/X _15010_/B1 vssd1 vssd1 vccd1 vccd1 _14990_/Y sky130_fd_sc_hd__a21oi_4
Xfanout1248 _08930_/Y vssd1 vssd1 vccd1 vccd1 _16820_/A3 sky130_fd_sc_hd__buf_4
XFILLER_259_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1259 _13807_/A vssd1 vssd1 vccd1 vccd1 _13937_/A sky130_fd_sc_hd__buf_4
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13941_ _13941_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _13941_/X sky130_fd_sc_hd__or2_1
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16660_ _19242_/Q _16664_/C vssd1 vssd1 vccd1 vccd1 _16662_/B sky130_fd_sc_hd__nor2_1
XFILLER_234_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13872_ _17916_/Q _13971_/A2 _13870_/Y _13871_/Y _13579_/A vssd1 vssd1 vccd1 vccd1
+ _13872_/X sky130_fd_sc_hd__a221o_4
XFILLER_90_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15611_ _15591_/A _15590_/B _15590_/A vssd1 vssd1 vccd1 vccd1 _15612_/B sky130_fd_sc_hd__o21ba_2
XFILLER_262_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12823_ _12823_/A _12823_/B vssd1 vssd1 vccd1 vccd1 _12823_/Y sky130_fd_sc_hd__nand2_1
XFILLER_222_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16591_ _17691_/A _16591_/B vssd1 vssd1 vccd1 vccd1 _16591_/Y sky130_fd_sc_hd__nand2_2
XFILLER_234_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18330_ _19609_/CLK _18330_/D vssd1 vssd1 vccd1 vccd1 _18330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _15540_/Y _15542_/B vssd1 vssd1 vccd1 vccd1 _15544_/A sky130_fd_sc_hd__nand2b_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12755_/A _12754_/B vssd1 vssd1 vccd1 vccd1 _12754_/Y sky130_fd_sc_hd__nand2_2
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11705_ _11704_/A _14345_/B vssd1 vssd1 vccd1 vccd1 _11705_/Y sky130_fd_sc_hd__nand2b_1
X_18261_ _19643_/CLK _18261_/D vssd1 vssd1 vccd1 vccd1 _18261_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12685_ _12675_/X _12684_/Y _13089_/A vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__mux2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15473_ _15445_/A _15445_/B _15444_/A vssd1 vssd1 vccd1 vccd1 _15474_/B sky130_fd_sc_hd__o21ai_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_144_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19492_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17212_ _19422_/Q fanout534/X _17547_/A _17212_/B2 vssd1 vssd1 vccd1 vccd1 _17213_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_11636_ _11636_/A _11636_/B vssd1 vssd1 vccd1 vccd1 _13860_/A sky130_fd_sc_hd__nand2_8
X_14424_ _14424_/A _17231_/A vssd1 vssd1 vccd1 vccd1 _18276_/D sky130_fd_sc_hd__nor2_4
X_18192_ _19608_/CLK _18192_/D vssd1 vssd1 vccd1 vccd1 _18192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17143_ _19399_/Q _17124_/B _17428_/A _17158_/B2 vssd1 vssd1 vccd1 vccd1 _17144_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_129_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14355_ _18207_/Q _16529_/A0 _14383_/S vssd1 vssd1 vccd1 vccd1 _18207_/D sky130_fd_sc_hd__mux2_1
X_11567_ _11565_/X _11566_/X _11567_/S vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__mux2_1
XFILLER_171_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13306_ _17835_/Q _13821_/B _13305_/X vssd1 vssd1 vccd1 vccd1 _13306_/X sky130_fd_sc_hd__o21a_1
XFILLER_183_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10518_ _12320_/B _10518_/B vssd1 vssd1 vccd1 vccd1 _10518_/Y sky130_fd_sc_hd__nor2_1
X_14286_ _11452_/B _18145_/Q _14304_/S vssd1 vssd1 vccd1 vccd1 _18145_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17074_ _17579_/A _17074_/A2 _17073_/X _17338_/A vssd1 vssd1 vccd1 vccd1 _19370_/D
+ sky130_fd_sc_hd__o211a_1
X_11498_ _11498_/A1 _18145_/Q _18791_/Q _09966_/S vssd1 vssd1 vccd1 vccd1 _11498_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16025_ _18734_/Q _18726_/Q _16034_/S vssd1 vssd1 vccd1 vccd1 _16025_/X sky130_fd_sc_hd__mux2_1
X_13237_ _15330_/A _13236_/A _13237_/B1 vssd1 vssd1 vccd1 vccd1 _13255_/A sky130_fd_sc_hd__o21ai_1
X_10449_ _11365_/B2 _10414_/A2 _10448_/X _11133_/B2 vssd1 vssd1 vccd1 vccd1 _13775_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13168_ _19530_/Q _13372_/S vssd1 vssd1 vccd1 vccd1 _13168_/X sky130_fd_sc_hd__or2_1
XFILLER_152_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12119_ _17833_/Q _12120_/C _17834_/Q vssd1 vssd1 vccd1 vccd1 _12121_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17976_ _18627_/CLK _17976_/D vssd1 vssd1 vccd1 vccd1 _17976_/Q sky130_fd_sc_hd__dfxtp_1
X_13099_ _09476_/X _13292_/A2 _13098_/X _13256_/B1 _17926_/Q vssd1 vssd1 vccd1 vccd1
+ _13100_/B sky130_fd_sc_hd__a32o_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1760 _17912_/Q vssd1 vssd1 vccd1 vccd1 _09099_/A sky130_fd_sc_hd__clkbuf_16
X_16927_ _19316_/Q _17181_/B _16927_/S vssd1 vssd1 vccd1 vccd1 _16928_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1771 _17909_/Q vssd1 vssd1 vccd1 vccd1 _10471_/S sky130_fd_sc_hd__buf_12
Xfanout1782 _12962_/A0 vssd1 vssd1 vccd1 vccd1 _10373_/S sky130_fd_sc_hd__buf_12
XFILLER_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1793 _17903_/Q vssd1 vssd1 vccd1 vccd1 _09494_/A sky130_fd_sc_hd__buf_12
X_19646_ _19646_/CLK _19646_/D vssd1 vssd1 vccd1 vccd1 _19646_/Q sky130_fd_sc_hd__dfxtp_1
X_16858_ _16967_/S _17565_/B vssd1 vssd1 vccd1 vccd1 _16858_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15809_ _18601_/Q _16500_/A0 _15829_/S vssd1 vssd1 vccd1 vccd1 _18601_/D sky130_fd_sc_hd__mux2_1
X_19577_ _19609_/CLK _19577_/D vssd1 vssd1 vccd1 vccd1 _19577_/Q sky130_fd_sc_hd__dfxtp_1
X_16789_ _19284_/Q _16791_/C _16788_/Y vssd1 vssd1 vccd1 vccd1 _19284_/D sky130_fd_sc_hd__a21oi_1
XFILLER_225_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09330_ _09908_/A1 _09652_/A _09329_/X _09908_/B1 _18381_/Q vssd1 vssd1 vccd1 vccd1
+ _09331_/B sky130_fd_sc_hd__o32a_1
X_18528_ _19231_/CLK _18528_/D vssd1 vssd1 vccd1 vccd1 _18528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09261_ _09254_/X _09260_/X _09251_/X _09257_/X _12466_/A0 _12408_/A vssd1 vssd1
+ vccd1 vccd1 _09261_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18459_ _19575_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09192_ _09643_/A _11812_/A _09191_/Y _09946_/B1 vssd1 vssd1 vccd1 vccd1 _12599_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08976_ _10427_/C1 _08975_/X _11417_/B1 vssd1 vssd1 vccd1 vccd1 _08977_/B sky130_fd_sc_hd__a21o_1
XFILLER_76_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _11172_/A1 _17764_/Q _09680_/B1 _18313_/Q vssd1 vssd1 vccd1 vccd1 _09528_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _11397_/A1 _09455_/X _09456_/X _09458_/X vssd1 vssd1 vccd1 vccd1 _09459_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12470_ _16852_/A _14675_/C _12468_/Y vssd1 vssd1 vccd1 vccd1 _12538_/A sky130_fd_sc_hd__o21ai_4
XFILLER_177_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11421_ _11498_/A1 _18146_/Q _18792_/Q _09966_/S vssd1 vssd1 vccd1 vccd1 _11421_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14140_ _17690_/A0 _18079_/Q _14140_/S vssd1 vssd1 vccd1 vccd1 _18079_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11352_ _11352_/A1 _18953_/Q _18218_/Q _11353_/B2 vssd1 vssd1 vccd1 vccd1 _11352_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10303_ _11495_/B1 _10285_/X _10286_/X _10296_/X _10302_/X vssd1 vssd1 vccd1 vccd1
+ _10303_/X sky130_fd_sc_hd__o32a_4
XFILLER_192_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14071_ _17688_/A0 _18013_/Q _14072_/S vssd1 vssd1 vccd1 vccd1 _18013_/D sky130_fd_sc_hd__mux2_1
X_11283_ _11284_/A1 _19633_/Q _18922_/Q _11284_/B2 vssd1 vssd1 vccd1 vccd1 _11283_/X
+ sky130_fd_sc_hd__a22o_1
X_13022_ _17860_/Q _13945_/A2 _13011_/X _13303_/B2 _13952_/B1 vssd1 vssd1 vccd1 vccd1
+ _13023_/B sky130_fd_sc_hd__a221o_1
XFILLER_3_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10234_ _11218_/A _10234_/B vssd1 vssd1 vccd1 vccd1 _10235_/B sky130_fd_sc_hd__nor2_1
XFILLER_267_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1001 _10414_/A2 vssd1 vssd1 vccd1 vccd1 _16618_/A0 sky130_fd_sc_hd__buf_2
XFILLER_3_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17830_ _19306_/CLK _17830_/D vssd1 vssd1 vccd1 vccd1 _17830_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1012 _15047_/Y vssd1 vssd1 vccd1 vccd1 _15070_/S sky130_fd_sc_hd__buf_4
X_10165_ _11064_/B1 _10163_/Y _10164_/X vssd1 vssd1 vccd1 vccd1 _10165_/X sky130_fd_sc_hd__o21a_1
XFILLER_117_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1023 _11558_/X vssd1 vssd1 vccd1 vccd1 _17690_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_239_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1034 _09611_/B vssd1 vssd1 vccd1 vccd1 _16465_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1045 _08958_/X vssd1 vssd1 vccd1 vccd1 _11133_/B2 sky130_fd_sc_hd__buf_8
Xfanout1056 _15523_/S vssd1 vssd1 vccd1 vccd1 _15716_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17761_ _19148_/CLK _17761_/D vssd1 vssd1 vccd1 vccd1 _17761_/Q sky130_fd_sc_hd__dfxtp_1
X_10096_ _10253_/A _10095_/X _10094_/X vssd1 vssd1 vccd1 vccd1 _10096_/Y sky130_fd_sc_hd__o21ai_1
X_14973_ _14973_/A1 _13856_/Y _14973_/B1 _18654_/Q _14973_/C1 vssd1 vssd1 vccd1 vccd1
+ _14973_/X sky130_fd_sc_hd__a221o_1
Xfanout1067 _12741_/Y vssd1 vssd1 vccd1 vccd1 _13486_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1078 _17659_/A0 vssd1 vssd1 vccd1 vccd1 _16526_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_281_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1089 _16595_/A0 vssd1 vssd1 vccd1 vccd1 _17695_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19500_ _19533_/CLK _19500_/D vssd1 vssd1 vccd1 vccd1 _19500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16712_ _19256_/Q _16717_/D _19257_/Q vssd1 vssd1 vccd1 vccd1 _16714_/B sky130_fd_sc_hd__a21oi_1
XFILLER_263_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13924_ _19486_/Q _12529_/Y _12578_/Y _19358_/Q _13923_/X vssd1 vssd1 vccd1 vccd1
+ _13924_/X sky130_fd_sc_hd__a221o_1
X_17692_ _17692_/A0 _19618_/Q _17723_/S vssd1 vssd1 vccd1 vccd1 _19618_/D sky130_fd_sc_hd__mux2_1
XFILLER_247_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19431_ _19530_/CLK _19431_/D vssd1 vssd1 vccd1 vccd1 _19431_/Q sky130_fd_sc_hd__dfxtp_1
X_16643_ _19237_/Q _19236_/Q _16643_/C vssd1 vssd1 vccd1 vccd1 _16649_/C sky130_fd_sc_hd__and3_1
X_13855_ _13928_/A1 _13844_/X _13846_/Y _13854_/Y vssd1 vssd1 vccd1 vccd1 _14030_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_207_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19362_ _19458_/CLK _19362_/D vssd1 vssd1 vccd1 vccd1 _19362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12806_ _12804_/X _12805_/X _12943_/S vssd1 vssd1 vccd1 vccd1 _12806_/X sky130_fd_sc_hd__mux2_1
XFILLER_250_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16574_ _16607_/A0 _19178_/Q _16585_/S vssd1 vssd1 vccd1 vccd1 _19178_/D sky130_fd_sc_hd__mux2_1
X_10998_ _18425_/Q _11479_/B _10997_/X _11002_/C1 vssd1 vssd1 vccd1 vccd1 _10998_/X
+ sky130_fd_sc_hd__o211a_1
X_13786_ _19322_/Q _13174_/A _13779_/X _13785_/X vssd1 vssd1 vccd1 vccd1 _13786_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_90_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18313_ _19201_/CLK _18313_/D vssd1 vssd1 vccd1 vccd1 _18313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _18580_/Q _15718_/A2 _15524_/X _17354_/A vssd1 vssd1 vccd1 vccd1 _18580_/D
+ sky130_fd_sc_hd__o211a_1
X_19293_ _19327_/CLK _19293_/D vssd1 vssd1 vccd1 vccd1 _19293_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12727_/X _12988_/B _13089_/A vssd1 vssd1 vccd1 vccd1 _12737_/X sky130_fd_sc_hd__mux2_2
XFILLER_124_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _19047_/CLK _18244_/D vssd1 vssd1 vccd1 vccd1 _18244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15456_ _15456_/A _15456_/B _15456_/C _15456_/D vssd1 vssd1 vccd1 vccd1 _15457_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_230_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12668_ _12599_/B _12640_/B _12729_/B vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14407_ _16614_/A0 _18258_/Q _14412_/S vssd1 vssd1 vccd1 vccd1 _18258_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18175_ _19203_/CLK _18175_/D vssd1 vssd1 vccd1 vccd1 _18175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11619_ _11282_/A _11617_/X _11618_/X _11285_/S vssd1 vssd1 vccd1 vccd1 _11619_/X
+ sky130_fd_sc_hd__a211o_1
X_15387_ _15387_/A _15387_/B vssd1 vssd1 vccd1 vccd1 _15456_/B sky130_fd_sc_hd__xnor2_1
XFILLER_129_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12599_ _12599_/A _12599_/B vssd1 vssd1 vccd1 vccd1 _12622_/A sky130_fd_sc_hd__nand2_1
XFILLER_117_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17126_ _17157_/A _17563_/A vssd1 vssd1 vccd1 vccd1 _17404_/A sky130_fd_sc_hd__nand2_1
XFILLER_274_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14338_ _18195_/Q _15832_/A1 _14338_/S vssd1 vssd1 vccd1 vccd1 _18195_/D sky130_fd_sc_hd__mux2_1
XFILLER_184_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17057_ _19362_/Q _17113_/B vssd1 vssd1 vccd1 vccd1 _17057_/X sky130_fd_sc_hd__or2_1
X_14269_ _18306_/Q _14268_/B _14268_/Y _17356_/A vssd1 vssd1 vccd1 vccd1 _18132_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16008_ _18719_/Q _15953_/B _16147_/A2 _18768_/Q _16018_/C1 vssd1 vssd1 vccd1 vccd1
+ _16008_/X sky130_fd_sc_hd__a221o_1
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19608_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08830_ _18503_/Q vssd1 vssd1 vccd1 vccd1 _08830_/Y sky130_fd_sc_hd__inv_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17959_ _17975_/CLK _17959_/D vssd1 vssd1 vccd1 vccd1 _17959_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1590 _11503_/S1 vssd1 vssd1 vccd1 vccd1 _11510_/S1 sky130_fd_sc_hd__buf_6
XFILLER_39_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19629_ _19629_/CLK _19629_/D vssd1 vssd1 vccd1 vccd1 _19629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09313_ _11518_/B2 _16204_/A0 _09312_/X _09523_/A vssd1 vssd1 vccd1 vccd1 _15284_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_179_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09244_ _18382_/Q _09908_/B1 _09243_/Y _09992_/A vssd1 vssd1 vccd1 vccd1 _09245_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_167_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09175_ _11017_/A1 _18604_/Q _18175_/Q _10099_/S vssd1 vssd1 vccd1 vccd1 _09175_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput104 dout0[7] vssd1 vssd1 vccd1 vccd1 input104/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput115 dout1[17] vssd1 vssd1 vccd1 vccd1 input115/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput126 dout1[27] vssd1 vssd1 vccd1 vccd1 input126/X sky130_fd_sc_hd__clkbuf_2
XFILLER_277_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput137 dout1[37] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_hd__buf_2
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput148 dout1[47] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_hd__buf_2
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput159 dout1[57] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_hd__buf_2
XFILLER_276_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08959_ _18543_/Q _18418_/Q _18027_/Q _17995_/Q _11503_/S0 _11510_/S1 vssd1 vssd1
+ vccd1 vccd1 _08959_/X sky130_fd_sc_hd__mux4_1
XFILLER_248_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _18741_/Q _11981_/B _16054_/A vssd1 vssd1 vccd1 vccd1 _16056_/B sky130_fd_sc_hd__and3_4
XFILLER_57_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10921_ _18551_/Q _11309_/S vssd1 vssd1 vccd1 vccd1 _10921_/X sky130_fd_sc_hd__or2_1
XFILLER_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13640_ _13968_/A1 _13622_/Y _13639_/X _13621_/X _13323_/B vssd1 vssd1 vccd1 vccd1
+ _13640_/X sky130_fd_sc_hd__a32o_2
X_10852_ _18459_/Q _18360_/Q _10853_/S vssd1 vssd1 vccd1 vccd1 _10852_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13571_ _12265_/B _13568_/A _13570_/X vssd1 vssd1 vccd1 vccd1 _13571_/Y sky130_fd_sc_hd__a21oi_1
X_10783_ _10850_/A1 _19152_/Q _11302_/S _19120_/Q vssd1 vssd1 vccd1 vccd1 _10783_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _15310_/A _15310_/B vssd1 vssd1 vccd1 vccd1 _15312_/B sky130_fd_sc_hd__nand2_1
XFILLER_188_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12522_ _08817_/Y _12851_/B _12576_/A _12577_/B _12577_/A vssd1 vssd1 vccd1 vccd1
+ _12522_/Y sky130_fd_sc_hd__a2111oi_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16621_/A0 _18904_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _18904_/D sky130_fd_sc_hd__mux2_1
XFILLER_169_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ _12318_/Y _15381_/A3 _08840_/Y vssd1 vssd1 vccd1 vccd1 _15243_/B sky130_fd_sc_hd__a21o_2
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12453_ _09494_/A _10061_/X _13446_/B vssd1 vssd1 vccd1 vccd1 _12453_/X sky130_fd_sc_hd__mux2_1
X_11404_ _11404_/A1 _18146_/Q _18792_/Q _11481_/C vssd1 vssd1 vccd1 vccd1 _11404_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12384_ _11695_/B _09652_/A _09002_/X _12432_/B1 _18388_/Q vssd1 vssd1 vccd1 vccd1
+ _12385_/C sky130_fd_sc_hd__o32a_1
XFILLER_166_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15172_ _17899_/Q _15328_/B _15328_/C _12761_/B _17912_/Q vssd1 vssd1 vccd1 vccd1
+ _15177_/A sky130_fd_sc_hd__a32o_2
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ _16540_/A0 _18062_/Q _14140_/S vssd1 vssd1 vccd1 vccd1 _18062_/D sky130_fd_sc_hd__mux2_1
X_11335_ _12756_/A _11337_/B _11489_/B1 _11334_/Y vssd1 vssd1 vccd1 vccd1 _12596_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18931_ _19641_/CLK _18931_/D vssd1 vssd1 vccd1 vccd1 _18931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14054_ _17671_/A0 _17996_/Q _14072_/S vssd1 vssd1 vccd1 vccd1 _17996_/D sky130_fd_sc_hd__mux2_1
X_11266_ _10745_/S _11265_/X _11279_/B1 vssd1 vssd1 vccd1 vccd1 _11266_/X sky130_fd_sc_hd__a21o_1
X_10217_ _18904_/Q _10217_/B vssd1 vssd1 vccd1 vccd1 _10217_/X sky130_fd_sc_hd__or2_1
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13005_ _14214_/A _09948_/B _12984_/X _13004_/Y _13292_/A2 vssd1 vssd1 vccd1 vccd1
+ _13005_/X sky130_fd_sc_hd__o221a_1
XFILLER_239_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18862_ _19632_/CLK _18862_/D vssd1 vssd1 vccd1 vccd1 _18862_/Q sky130_fd_sc_hd__dfxtp_1
X_11197_ _11277_/A1 _18149_/Q _18795_/Q _10717_/S vssd1 vssd1 vccd1 vccd1 _11197_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_279_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17813_ _19492_/CLK _17813_/D vssd1 vssd1 vccd1 vccd1 _17813_/Q sky130_fd_sc_hd__dfxtp_4
X_10148_ _10297_/A1 _10138_/X _10139_/X vssd1 vssd1 vccd1 vccd1 _10148_/X sky130_fd_sc_hd__o21a_1
XFILLER_255_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18793_ _19216_/CLK _18793_/D vssd1 vssd1 vccd1 vccd1 _18793_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17744_ _18644_/Q vssd1 vssd1 vccd1 vccd1 _18644_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_248_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14956_ _15006_/A1 _14955_/X _11715_/B vssd1 vssd1 vccd1 vccd1 _14956_/Y sky130_fd_sc_hd__o21ai_2
X_10079_ _13225_/A _11753_/B _13230_/S vssd1 vssd1 vccd1 vccd1 _10080_/B sky130_fd_sc_hd__o21ba_4
XFILLER_254_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13907_ _13891_/A _13860_/A _13860_/B _12659_/Y vssd1 vssd1 vccd1 vccd1 _13908_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_223_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17675_ _17708_/A0 _19602_/Q _17681_/S vssd1 vssd1 vccd1 vccd1 _19602_/D sky130_fd_sc_hd__mux2_1
X_14887_ _14887_/A vssd1 vssd1 vccd1 vccd1 _14887_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_250_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19414_ _19546_/CLK _19414_/D vssd1 vssd1 vccd1 vccd1 _19414_/Q sky130_fd_sc_hd__dfxtp_2
X_16626_ _19229_/Q input249/X _16627_/S vssd1 vssd1 vccd1 vccd1 _19229_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13838_ _13900_/C _13838_/B vssd1 vssd1 vccd1 vccd1 _13838_/X sky130_fd_sc_hd__or2_1
XFILLER_262_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19345_ _19507_/CLK _19345_/D vssd1 vssd1 vccd1 vccd1 _19345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16557_ _16557_/A0 _19162_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _19162_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13769_ _13323_/B _13768_/X _13760_/X vssd1 vssd1 vccd1 vccd1 _13769_/X sky130_fd_sc_hd__a21o_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15508_ _15487_/A _15508_/B vssd1 vssd1 vccd1 vccd1 _15508_/X sky130_fd_sc_hd__and2b_1
X_19276_ _19276_/CLK _19276_/D vssd1 vssd1 vccd1 vccd1 _19276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16488_ _16488_/A0 _19095_/Q _16488_/S vssd1 vssd1 vccd1 vccd1 _19095_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18227_ _19155_/CLK _18227_/D vssd1 vssd1 vccd1 vccd1 _18227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15439_ _15124_/B _15435_/X _15437_/X _15438_/Y vssd1 vssd1 vccd1 vccd1 _15439_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_129_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18158_ _19642_/CLK _18158_/D vssd1 vssd1 vccd1 vccd1 _18158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17109_ _19388_/Q _17115_/B vssd1 vssd1 vccd1 vccd1 _17109_/X sky130_fd_sc_hd__or2_1
XFILLER_190_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18089_ _18776_/CLK _18089_/D vssd1 vssd1 vccd1 vccd1 _18089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _09929_/X _09930_/X _08843_/A vssd1 vssd1 vccd1 vccd1 _09931_/X sky130_fd_sc_hd__a21o_1
XFILLER_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout805 _15817_/S vssd1 vssd1 vccd1 vccd1 _15833_/S sky130_fd_sc_hd__buf_12
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout816 _14351_/Y vssd1 vssd1 vccd1 vccd1 _14380_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_98_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _15120_/A _11788_/B _09861_/Y _10027_/B vssd1 vssd1 vccd1 vccd1 _09862_/X
+ sky130_fd_sc_hd__a211o_4
Xfanout827 _11990_/Y vssd1 vssd1 vccd1 vccd1 _12013_/S sky130_fd_sc_hd__clkbuf_8
Xfanout838 _17710_/A0 vssd1 vssd1 vccd1 vccd1 _17677_/A0 sky130_fd_sc_hd__clkbuf_4
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout849 _10837_/X vssd1 vssd1 vccd1 vccd1 _14510_/A0 sky130_fd_sc_hd__buf_4
XFILLER_285_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _19621_/Q _18910_/Q _09797_/S vssd1 vssd1 vccd1 vccd1 _09793_/X sky130_fd_sc_hd__mux2_1
XFILLER_274_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _18564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09227_ _09946_/B1 _15303_/A _09193_/X vssd1 vssd1 vccd1 vccd1 _09229_/B sky130_fd_sc_hd__o21ai_4
XFILLER_194_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09158_ _17962_/Q _11295_/A2 _08947_/A _17930_/Q _08946_/B vssd1 vssd1 vccd1 vccd1
+ _09158_/X sky130_fd_sc_hd__a221o_1
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09089_ _12408_/A _09285_/C vssd1 vssd1 vccd1 vccd1 _09089_/Y sky130_fd_sc_hd__nand2_8
XFILLER_218_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11120_ _11118_/X _11119_/X _11127_/S vssd1 vssd1 vccd1 vccd1 _11120_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _11511_/A _11046_/X _11050_/X vssd1 vssd1 vccd1 vccd1 _11053_/C sky130_fd_sc_hd__a21oi_1
XFILLER_150_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10002_ _10027_/A _19067_/Q _18971_/Q _11224_/B _11569_/S1 vssd1 vssd1 vccd1 vccd1
+ _10002_/X sky130_fd_sc_hd__o221a_1
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _17802_/Q _14809_/X _14993_/S vssd1 vssd1 vccd1 vccd1 _14810_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _18593_/Q _15791_/B vssd1 vssd1 vccd1 vccd1 _15790_/X sky130_fd_sc_hd__or2_1
XFILLER_190_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _14741_/A _14741_/B vssd1 vssd1 vccd1 vccd1 _14741_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _19227_/Q _11953_/A2 _14342_/C _11953_/B2 vssd1 vssd1 vccd1 vccd1 _11953_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ _13581_/A vssd1 vssd1 vccd1 vccd1 _10904_/Y sky130_fd_sc_hd__inv_2
X_17460_ _13402_/B _15118_/A _15117_/A _12053_/A _15116_/B vssd1 vssd1 vccd1 vccd1
+ _17460_/X sky130_fd_sc_hd__a221o_1
XFILLER_264_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _14688_/B _14680_/B _14672_/C _14681_/B vssd1 vssd1 vccd1 vccd1 _14672_/X
+ sky130_fd_sc_hd__and4bb_1
X_11884_ _11812_/X _11875_/A _11901_/B _11845_/X vssd1 vssd1 vccd1 vccd1 _11884_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16411_ _16609_/A0 _19020_/Q _16420_/S vssd1 vssd1 vccd1 vccd1 _19020_/D sky130_fd_sc_hd__mux2_1
XFILLER_233_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13623_ _13623_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13638_/B sky130_fd_sc_hd__or2_1
XFILLER_232_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10835_ _17972_/Q _11216_/A2 _11216_/B1 vssd1 vssd1 vccd1 vccd1 _10835_/X sky130_fd_sc_hd__a21o_1
X_17391_ _11824_/A _15118_/A _15117_/A _17790_/Q vssd1 vssd1 vccd1 vccd1 _17391_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19130_ _19163_/CLK _19130_/D vssd1 vssd1 vccd1 vccd1 _19130_/Q sky130_fd_sc_hd__dfxtp_1
X_16342_ _18954_/Q _17674_/A0 _16352_/S vssd1 vssd1 vccd1 vccd1 _18954_/D sky130_fd_sc_hd__mux2_1
XFILLER_198_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13554_ _19509_/Q _13947_/A2 _13947_/B1 _13553_/X vssd1 vssd1 vccd1 vccd1 _13554_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10766_ _11327_/S _10765_/X _10764_/X vssd1 vssd1 vccd1 vccd1 _10766_/X sky130_fd_sc_hd__o21a_1
XFILLER_186_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12505_ _13167_/A _13165_/B vssd1 vssd1 vccd1 vccd1 _12505_/Y sky130_fd_sc_hd__nor2_4
X_19061_ _19219_/CLK _19061_/D vssd1 vssd1 vccd1 vccd1 _19061_/Q sky130_fd_sc_hd__dfxtp_1
X_16273_ _11452_/B _18887_/Q _16288_/S vssd1 vssd1 vccd1 vccd1 _18887_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10697_ _10689_/S _10692_/X _10696_/X _09350_/S vssd1 vssd1 vccd1 vccd1 _10697_/X
+ sky130_fd_sc_hd__o211a_1
X_13485_ _13485_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _14146_/B sky130_fd_sc_hd__xnor2_1
XFILLER_201_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18012_ _19614_/CLK _18012_/D vssd1 vssd1 vccd1 vccd1 _18012_/Q sky130_fd_sc_hd__dfxtp_1
X_15224_ _18568_/Q _18567_/Q _15224_/C vssd1 vssd1 vccd1 vccd1 _15270_/C sky130_fd_sc_hd__and3_1
XFILLER_218_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12436_ _12437_/A _12587_/B vssd1 vssd1 vccd1 vccd1 _12436_/X sky130_fd_sc_hd__and2_1
XFILLER_126_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput408 _11984_/X vssd1 vssd1 vccd1 vccd1 jtag_tdo sky130_fd_sc_hd__buf_4
X_15155_ _15155_/A _15155_/B vssd1 vssd1 vccd1 vccd1 _15156_/B sky130_fd_sc_hd__nand2_1
Xoutput419 _18489_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[18] sky130_fd_sc_hd__buf_4
X_12367_ _12408_/B _12367_/B vssd1 vssd1 vccd1 vccd1 _12367_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14106_ _17722_/A0 _18046_/Q _14106_/S vssd1 vssd1 vccd1 vccd1 _18046_/D sky130_fd_sc_hd__mux2_1
X_11318_ _11327_/S _19177_/Q _11325_/S vssd1 vssd1 vccd1 vccd1 _11318_/X sky130_fd_sc_hd__and3_1
X_12298_ _18083_/Q _12277_/B _14934_/C _18506_/Q vssd1 vssd1 vccd1 vccd1 _14675_/C
+ sky130_fd_sc_hd__a22o_4
X_15086_ _19381_/Q _15086_/B _15086_/C vssd1 vssd1 vccd1 vccd1 _15086_/X sky130_fd_sc_hd__and3_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18914_ _19625_/CLK _18914_/D vssd1 vssd1 vccd1 vccd1 _18914_/Q sky130_fd_sc_hd__dfxtp_1
X_14037_ _17983_/Q _14020_/B _14036_/Y _14037_/C1 vssd1 vssd1 vccd1 vccd1 _17983_/D
+ sky130_fd_sc_hd__o211a_1
X_11249_ _18858_/Q _18890_/Q _11249_/S vssd1 vssd1 vccd1 vccd1 _11249_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18845_ _19588_/CLK _18845_/D vssd1 vssd1 vccd1 vccd1 _18845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18776_ _18776_/CLK _18776_/D vssd1 vssd1 vccd1 vccd1 _18776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_282_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15988_ _18709_/Q _16016_/A2 _16004_/B1 _18758_/Q _16004_/C1 vssd1 vssd1 vccd1 vccd1
+ _15988_/X sky130_fd_sc_hd__a221o_1
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17727_ _18627_/Q vssd1 vssd1 vccd1 vccd1 _18627_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_282_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14939_ _14979_/A1 _18272_/Q _14938_/Y _11712_/A vssd1 vssd1 vccd1 vccd1 _14939_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_264_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17658_ _17658_/A _17691_/A vssd1 vssd1 vccd1 vccd1 _17658_/Y sky130_fd_sc_hd__nand2_8
XFILLER_251_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16609_ _16609_/A0 _19212_/Q _16618_/S vssd1 vssd1 vccd1 vccd1 _19212_/D sky130_fd_sc_hd__mux2_1
XFILLER_196_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17589_ _17589_/A _17589_/B vssd1 vssd1 vccd1 vccd1 _17589_/X sky130_fd_sc_hd__or2_1
X_19328_ _19458_/CLK _19328_/D vssd1 vssd1 vccd1 vccd1 _19328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_259_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19259_ _19261_/CLK _19259_/D vssd1 vssd1 vccd1 vccd1 _19259_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_176_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09012_ _09012_/A _09991_/A _09012_/C vssd1 vssd1 vccd1 vccd1 _09012_/X sky130_fd_sc_hd__or3_1
XFILLER_117_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09914_ _09935_/A _09912_/X _09913_/X _09914_/C1 vssd1 vssd1 vccd1 vccd1 _09914_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout602 _11696_/X vssd1 vssd1 vccd1 vccd1 _17724_/B sky130_fd_sc_hd__buf_8
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout613 _11654_/Y vssd1 vssd1 vccd1 vccd1 _11799_/A sky130_fd_sc_hd__buf_8
XFILLER_120_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout624 _17008_/A2 vssd1 vssd1 vccd1 vccd1 _17044_/A2 sky130_fd_sc_hd__buf_4
XFILLER_259_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout635 _11652_/Y vssd1 vssd1 vccd1 vccd1 _11826_/A sky130_fd_sc_hd__buf_6
XFILLER_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout646 _17107_/B vssd1 vssd1 vccd1 vccd1 _17115_/B sky130_fd_sc_hd__buf_4
XFILLER_219_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout657 _12580_/Y vssd1 vssd1 vccd1 vccd1 _13277_/S sky130_fd_sc_hd__buf_4
X_09845_ _09842_/X _09844_/X _09845_/S vssd1 vssd1 vccd1 vccd1 _09845_/X sky130_fd_sc_hd__mux2_1
Xfanout668 _11859_/A vssd1 vssd1 vccd1 vccd1 _11865_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout679 _13951_/A2 vssd1 vssd1 vccd1 vccd1 _13884_/A2 sky130_fd_sc_hd__buf_8
XFILLER_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09776_ _08852_/Y _11706_/C _10027_/B _09775_/X vssd1 vssd1 vccd1 vccd1 _09776_/X
+ sky130_fd_sc_hd__a211o_2
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10620_ _11584_/A1 _18156_/Q _18802_/Q _10619_/S vssd1 vssd1 vccd1 vccd1 _10620_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10551_ _11312_/A1 _17782_/Q _09108_/B _18331_/Q vssd1 vssd1 vccd1 vccd1 _10551_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13270_ _12440_/X _13265_/Y _13269_/X vssd1 vssd1 vccd1 vccd1 _13270_/X sky130_fd_sc_hd__a21bo_1
X_10482_ _10480_/X _10481_/X _10632_/S vssd1 vssd1 vccd1 vccd1 _10483_/B sky130_fd_sc_hd__mux2_1
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12221_ _17872_/Q _12224_/C _12241_/A vssd1 vssd1 vccd1 vccd1 _12221_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ _17845_/Q _17846_/Q _12152_/C vssd1 vssd1 vccd1 vccd1 _12154_/B sky130_fd_sc_hd__and3_2
XFILLER_2_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_169_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19484_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11103_ _11103_/A _11841_/A vssd1 vssd1 vccd1 vccd1 _11103_/Y sky130_fd_sc_hd__nor2_1
X_16960_ _16960_/A _16960_/B vssd1 vssd1 vccd1 vccd1 _19324_/D sky130_fd_sc_hd__and2_1
X_12083_ _17819_/Q _12087_/B vssd1 vssd1 vccd1 vccd1 _12083_/X sky130_fd_sc_hd__or2_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15911_ _15911_/A _15947_/S _15923_/C vssd1 vssd1 vccd1 vccd1 _15911_/X sky130_fd_sc_hd__and3_1
X_11034_ _11511_/A _11034_/B vssd1 vssd1 vccd1 vccd1 _11039_/A sky130_fd_sc_hd__and2_1
XFILLER_238_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16891_ _19307_/Q _17581_/A _16971_/S vssd1 vssd1 vccd1 vccd1 _16892_/B sky130_fd_sc_hd__mux2_1
XFILLER_238_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18630_ _19147_/CLK _18630_/D vssd1 vssd1 vccd1 vccd1 _18630_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _18742_/Q _12276_/A _16877_/B1 input215/X vssd1 vssd1 vccd1 vccd1 _15843_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_264_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18561_ _19615_/CLK _18561_/D vssd1 vssd1 vccd1 vccd1 _18561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_252_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _15789_/B1 _15791_/B _15772_/X _15751_/A vssd1 vssd1 vccd1 vccd1 _15773_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12985_ _12985_/A _12985_/B vssd1 vssd1 vccd1 vccd1 _14142_/A sky130_fd_sc_hd__xnor2_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17512_ _18125_/Q _17545_/C1 _17510_/X _17511_/X vssd1 vssd1 vccd1 vccd1 _17512_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_233_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _18104_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14724_/X sky130_fd_sc_hd__or2_1
X_18492_ _19286_/CLK _18492_/D vssd1 vssd1 vccd1 vccd1 _18492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _11953_/B2 _11840_/B _11953_/A2 input222/X vssd1 vssd1 vccd1 vccd1 _11936_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_220_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_540 _11940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _17443_/A _17453_/B vssd1 vssd1 vccd1 vccd1 _17443_/Y sky130_fd_sc_hd__nand2_1
XFILLER_221_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14655_ _17714_/A0 _18461_/Q _14660_/S vssd1 vssd1 vccd1 vccd1 _18461_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _11952_/A2 _11901_/A _11866_/X vssd1 vssd1 vccd1 vccd1 _11868_/B sky130_fd_sc_hd__a21oi_4
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ _18121_/Q _18120_/Q _13606_/C vssd1 vssd1 vccd1 vccd1 _13642_/B sky130_fd_sc_hd__and3_1
X_17374_ _17374_/A _17374_/B vssd1 vssd1 vccd1 vccd1 _19484_/D sky130_fd_sc_hd__and2_1
X_10818_ _10815_/X _10816_/X _10817_/X _10663_/S _11607_/S vssd1 vssd1 vccd1 vccd1
+ _10818_/X sky130_fd_sc_hd__a221o_1
XFILLER_159_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14586_ _14586_/A _14586_/B vssd1 vssd1 vccd1 vccd1 _18401_/D sky130_fd_sc_hd__or2_1
X_11798_ _11816_/A _11798_/B vssd1 vssd1 vccd1 vccd1 _11865_/B sky130_fd_sc_hd__nor2_8
XFILLER_201_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19113_ _19600_/CLK _19113_/D vssd1 vssd1 vccd1 vccd1 _19113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16325_ _17723_/A0 _18938_/Q _16325_/S vssd1 vssd1 vccd1 vccd1 _18938_/D sky130_fd_sc_hd__mux2_1
X_13537_ _13602_/B2 _13353_/X _13356_/X _12835_/A _13536_/X vssd1 vssd1 vccd1 vccd1
+ _13537_/X sky130_fd_sc_hd__o221a_1
X_10749_ _11210_/A1 _10713_/A2 _10748_/Y _11055_/B2 vssd1 vssd1 vccd1 vccd1 _13647_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19044_ _19208_/CLK _19044_/D vssd1 vssd1 vccd1 vccd1 _19044_/Q sky130_fd_sc_hd__dfxtp_1
X_16256_ _16455_/A1 _18871_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _18871_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13468_ _14155_/B _12756_/Y _13468_/S vssd1 vssd1 vccd1 vccd1 _13468_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15207_ _15207_/A _15207_/B vssd1 vssd1 vccd1 vccd1 _15207_/Y sky130_fd_sc_hd__xnor2_1
X_12419_ _17914_/Q _12427_/A _12418_/Y _12428_/C1 vssd1 vssd1 vccd1 vccd1 _17914_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16187_ _16617_/A0 _18804_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _18804_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13399_ _13406_/B _13399_/B vssd1 vssd1 vccd1 vccd1 _13399_/X sky130_fd_sc_hd__or2_1
XFILLER_126_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15138_ _15307_/B _15138_/B _15138_/C vssd1 vssd1 vccd1 vccd1 _15138_/X sky130_fd_sc_hd__or3_1
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15069_ _18553_/Q _17680_/A0 _15079_/S vssd1 vssd1 vccd1 vccd1 _18553_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09630_ _09690_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09630_/Y sky130_fd_sc_hd__nor2_1
X_18828_ _19637_/CLK _18828_/D vssd1 vssd1 vccd1 vccd1 _18828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09561_ _12613_/B _09561_/B vssd1 vssd1 vccd1 vccd1 _11742_/B sky130_fd_sc_hd__or2_2
X_18759_ _18761_/CLK _18759_/D vssd1 vssd1 vccd1 vccd1 _18759_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_283_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09492_ _19041_/Q _19009_/Q _09952_/S vssd1 vssd1 vccd1 vccd1 _09492_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1408 fanout1415/X vssd1 vssd1 vccd1 vccd1 _10176_/S sky130_fd_sc_hd__buf_6
XFILLER_259_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1419 _11403_/S vssd1 vssd1 vccd1 vccd1 _09252_/S sky130_fd_sc_hd__buf_4
XFILLER_59_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09828_ _11566_/A1 _19620_/Q _18909_/Q _10001_/S vssd1 vssd1 vccd1 vccd1 _09829_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout498 _11949_/B1 vssd1 vssd1 vccd1 vccd1 _11953_/A2 sky130_fd_sc_hd__buf_6
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09759_ _11568_/A _09758_/X _11563_/B1 vssd1 vssd1 vccd1 vccd1 _09759_/X sky130_fd_sc_hd__o21a_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12770_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__and2_1
XFILLER_243_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11704_/A _11968_/B2 _11720_/X _18515_/Q vssd1 vssd1 vccd1 vccd1 _11721_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14440_ _18579_/Q _14452_/B vssd1 vssd1 vccd1 vccd1 _18292_/D sky130_fd_sc_hd__and2_1
XFILLER_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11653_/A _11653_/B vssd1 vssd1 vccd1 vccd1 _11652_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10603_ _10603_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _13727_/A sky130_fd_sc_hd__nor2_8
XFILLER_11_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14371_ _18223_/Q _17711_/A0 _14383_/S vssd1 vssd1 vccd1 vccd1 _18223_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11583_ _11583_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16110_ _16078_/X _16109_/Y _16110_/B1 vssd1 vssd1 vccd1 vccd1 _18757_/D sky130_fd_sc_hd__a21oi_1
X_13322_ _15426_/B _13323_/B vssd1 vssd1 vccd1 vccd1 _13322_/Y sky130_fd_sc_hd__nor2_4
X_10534_ _19642_/Q _18931_/Q _10619_/S vssd1 vssd1 vccd1 vccd1 _10534_/X sky130_fd_sc_hd__mux2_1
X_17090_ _17175_/B _17116_/A2 _17089_/X _17354_/A vssd1 vssd1 vccd1 vccd1 _19378_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16041_ _16041_/A _16063_/B vssd1 vssd1 vccd1 vccd1 _16041_/X sky130_fd_sc_hd__or2_1
XFILLER_109_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10465_ _10471_/S _10463_/X _10464_/X vssd1 vssd1 vccd1 vccd1 _10465_/X sky130_fd_sc_hd__o21a_1
X_13253_ _12587_/Y _13238_/X _13253_/B1 vssd1 vssd1 vccd1 vccd1 _13253_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12204_ _17865_/Q _12202_/B _12203_/Y vssd1 vssd1 vccd1 vccd1 _17865_/D sky130_fd_sc_hd__o21a_1
XFILLER_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10396_ _11312_/A1 _18159_/Q _18805_/Q _10864_/S vssd1 vssd1 vccd1 vccd1 _10396_/X
+ sky130_fd_sc_hd__a22o_1
X_13184_ _13079_/A _13182_/Y _13183_/X _13147_/A _13254_/B2 vssd1 vssd1 vccd1 vccd1
+ _13185_/D sky130_fd_sc_hd__a32o_1
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ _17839_/Q _12136_/C _17840_/Q vssd1 vssd1 vccd1 vccd1 _12137_/B sky130_fd_sc_hd__a21oi_1
XFILLER_2_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17992_ _19213_/CLK _17992_/D vssd1 vssd1 vccd1 vccd1 _17992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16943_ _19320_/Q _17193_/B _16947_/S vssd1 vssd1 vccd1 vccd1 _16944_/B sky130_fd_sc_hd__mux2_1
XFILLER_278_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12066_ _09457_/B _12088_/A2 _12065_/X _17328_/A vssd1 vssd1 vccd1 vccd1 _17810_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11017_ _11017_/A1 _18151_/Q _18797_/Q _11481_/C vssd1 vssd1 vccd1 vccd1 _11017_/X
+ sky130_fd_sc_hd__a22o_1
X_16874_ _16848_/S _17927_/Q _16873_/X vssd1 vssd1 vccd1 vccd1 _17573_/A sky130_fd_sc_hd__o21a_4
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15825_ _18617_/Q _17715_/A0 _15833_/S vssd1 vssd1 vccd1 vccd1 _18617_/D sky130_fd_sc_hd__mux2_1
X_18613_ _18613_/CLK _18613_/D vssd1 vssd1 vccd1 vccd1 _18613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19593_ _19614_/CLK _19593_/D vssd1 vssd1 vccd1 vccd1 _19593_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18544_ _19565_/CLK _18544_/D vssd1 vssd1 vccd1 vccd1 _18544_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _15756_/A _15756_/B vssd1 vssd1 vccd1 vccd1 _15757_/B sky130_fd_sc_hd__nand2_1
XFILLER_280_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ _19526_/Q _13372_/S vssd1 vssd1 vccd1 vccd1 _12968_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_66_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19636_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14707_ input54/X input69/X _14784_/S vssd1 vssd1 vccd1 vccd1 _14708_/B sky130_fd_sc_hd__mux2_8
X_18475_ _19319_/CLK _18475_/D vssd1 vssd1 vccd1 vccd1 _18475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11919_ _14667_/A1 _11919_/B _15835_/A vssd1 vssd1 vccd1 vccd1 _11919_/X sky130_fd_sc_hd__and3b_1
XFILLER_206_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15687_ _15687_/A _15687_/B vssd1 vssd1 vccd1 vccd1 _15725_/B sky130_fd_sc_hd__or2_1
XFILLER_61_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_370 _18203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12899_ _14153_/A _12899_/B _12898_/X vssd1 vssd1 vccd1 vccd1 _12899_/X sky130_fd_sc_hd__or3b_2
XANTENNA_381 _15010_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_392 _09004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17426_ _18569_/Q _17461_/A2 _17426_/B1 vssd1 vssd1 vccd1 vccd1 _17426_/X sky130_fd_sc_hd__o21a_1
X_14638_ _17697_/A0 _18444_/Q _14660_/S vssd1 vssd1 vccd1 vccd1 _18444_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17357_ _19476_/Q _17181_/B _17379_/S vssd1 vssd1 vccd1 vccd1 _17358_/B sky130_fd_sc_hd__mux2_1
X_14569_ _18393_/Q _14575_/A2 _14575_/B1 input22/X vssd1 vssd1 vccd1 vccd1 _14570_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ _17706_/A0 _18921_/Q _16320_/S vssd1 vssd1 vccd1 vccd1 _18921_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17288_ _17286_/Y _17287_/X _17198_/A vssd1 vssd1 vccd1 vccd1 _19446_/D sky130_fd_sc_hd__a21oi_1
XFILLER_173_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19027_ _19219_/CLK _19027_/D vssd1 vssd1 vccd1 vccd1 _19027_/Q sky130_fd_sc_hd__dfxtp_1
X_16239_ _09105_/A _18854_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _18854_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _11556_/A _08990_/X _08991_/X _08940_/B _08929_/B vssd1 vssd1 vccd1 vccd1
+ _08992_/Y sky130_fd_sc_hd__a2111oi_4
XFILLER_130_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09613_ _10323_/A1 _19559_/Q _09688_/S _19591_/Q vssd1 vssd1 vccd1 vccd1 _09613_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _09553_/A _09544_/B vssd1 vssd1 vccd1 vccd1 _09544_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09475_ _12612_/B _09475_/B vssd1 vssd1 vccd1 vccd1 _11745_/B sky130_fd_sc_hd__nor2_4
XPHY_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10250_ _10248_/X _10249_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _10250_/X sky130_fd_sc_hd__mux2_2
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10181_ _18561_/Q _18436_/Q _18045_/Q _18013_/Q _10090_/S _11001_/C1 vssd1 vssd1
+ vccd1 vccd1 _10181_/X sky130_fd_sc_hd__mux4_1
XFILLER_278_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1205 _12753_/X vssd1 vssd1 vccd1 vccd1 _13912_/B1 sky130_fd_sc_hd__buf_8
XFILLER_132_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1216 _12442_/D vssd1 vssd1 vccd1 vccd1 _13863_/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout1227 _15481_/B vssd1 vssd1 vccd1 vccd1 _15112_/A sky130_fd_sc_hd__buf_4
Xfanout1238 _09899_/X vssd1 vssd1 vccd1 vccd1 _11216_/B1 sky130_fd_sc_hd__buf_4
Xfanout1249 _08930_/Y vssd1 vssd1 vccd1 vccd1 _11295_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13940_ _17950_/Q _13940_/A2 _13939_/X _14029_/C1 vssd1 vssd1 vccd1 vccd1 _17950_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13871_ _13938_/A _17531_/A vssd1 vssd1 vccd1 vccd1 _13871_/Y sky130_fd_sc_hd__nand2_1
XFILLER_235_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15610_ _15610_/A _15610_/B vssd1 vssd1 vccd1 vccd1 _15612_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12822_ _12821_/A _12721_/X _12821_/Y vssd1 vssd1 vccd1 vccd1 _12822_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16590_ _17723_/A0 _19194_/Q _16590_/S vssd1 vssd1 vccd1 vccd1 _19194_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15541_ _19475_/Q _19409_/Q vssd1 vssd1 vccd1 vccd1 _15542_/B sky130_fd_sc_hd__nand2_1
XFILLER_199_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12753_ _12755_/A _12754_/B vssd1 vssd1 vccd1 vccd1 _12753_/X sky130_fd_sc_hd__and2_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11704_ _11704_/A _14345_/B vssd1 vssd1 vccd1 vccd1 _14487_/B sky130_fd_sc_hd__nand2_1
X_18260_ _19641_/CLK _18260_/D vssd1 vssd1 vccd1 vccd1 _18260_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15472_ _15472_/A _15472_/B vssd1 vssd1 vccd1 vccd1 _15474_/A sky130_fd_sc_hd__nand2_1
XFILLER_199_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12684_ _12933_/A _12678_/X _12683_/X vssd1 vssd1 vccd1 vccd1 _12684_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_187_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17211_ _17211_/A _17211_/B vssd1 vssd1 vccd1 vccd1 _17547_/A sky130_fd_sc_hd__nand2_1
X_14423_ _14423_/A _14423_/B vssd1 vssd1 vccd1 vccd1 _18275_/D sky130_fd_sc_hd__nor2_4
X_18191_ _19644_/CLK _18191_/D vssd1 vssd1 vccd1 vccd1 _18191_/Q sky130_fd_sc_hd__dfxtp_1
X_11635_ _11635_/A _13891_/A vssd1 vssd1 vccd1 vccd1 _13904_/B sky130_fd_sc_hd__xnor2_4
XFILLER_168_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17142_ _17151_/A _17573_/A vssd1 vssd1 vccd1 vccd1 _17428_/A sky130_fd_sc_hd__nand2_2
X_14354_ _18206_/Q _17661_/A0 _14377_/S vssd1 vssd1 vccd1 vccd1 _18206_/D sky130_fd_sc_hd__mux2_1
XFILLER_196_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ _11566_/A1 _19162_/Q _11226_/S _19130_/Q vssd1 vssd1 vccd1 vccd1 _11566_/X
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_184_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17930_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13305_ _17867_/Q _13847_/A2 _13854_/B1 _13304_/X vssd1 vssd1 vccd1 vccd1 _13305_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10517_ _10515_/X _10516_/X _10668_/S vssd1 vssd1 vccd1 vccd1 _10518_/B sky130_fd_sc_hd__mux2_1
X_17073_ _19370_/Q _17073_/B vssd1 vssd1 vccd1 vccd1 _17073_/X sky130_fd_sc_hd__or2_1
X_14285_ _09105_/A _18144_/Q _14304_/S vssd1 vssd1 vccd1 vccd1 _18144_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11497_ _11497_/A1 _19207_/Q _19175_/Q _09973_/S vssd1 vssd1 vccd1 vccd1 _11497_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_113_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18501_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16024_ _16020_/A _16056_/B _18727_/Q vssd1 vssd1 vccd1 vccd1 _16024_/X sky130_fd_sc_hd__a21o_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13236_ _13236_/A vssd1 vssd1 vccd1 vccd1 _13236_/Y sky130_fd_sc_hd__inv_2
X_10448_ _11279_/B1 _10431_/X _10446_/X _10447_/Y vssd1 vssd1 vccd1 vccd1 _10448_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13167_ _13167_/A _13167_/B vssd1 vssd1 vccd1 vccd1 _13174_/B sky130_fd_sc_hd__nor2_1
XFILLER_269_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10379_ _10381_/A _12653_/B vssd1 vssd1 vccd1 vccd1 _11550_/A sky130_fd_sc_hd__nor2_4
XFILLER_285_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ _17833_/Q _12120_/C _12117_/Y vssd1 vssd1 vccd1 vccd1 _17833_/D sky130_fd_sc_hd__o21a_1
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17975_ _17975_/CLK _17975_/D vssd1 vssd1 vccd1 vccd1 _17975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13098_ _12447_/Y _13085_/X _13097_/X _13080_/X vssd1 vssd1 vccd1 vccd1 _13098_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_242_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1750 _17920_/Q vssd1 vssd1 vccd1 vccd1 _09031_/S sky130_fd_sc_hd__buf_8
XFILLER_66_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16926_ _16848_/S _17940_/Q _16925_/X vssd1 vssd1 vccd1 vccd1 _17181_/B sky130_fd_sc_hd__o21a_4
X_12049_ _17802_/Q _12073_/B vssd1 vssd1 vccd1 vccd1 _12049_/X sky130_fd_sc_hd__or2_1
Xfanout1761 _09777_/A vssd1 vssd1 vccd1 vccd1 _12408_/A sky130_fd_sc_hd__buf_12
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1772 _12471_/A0 vssd1 vssd1 vccd1 vccd1 _11173_/S sky130_fd_sc_hd__buf_8
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1783 _17907_/Q vssd1 vssd1 vccd1 vccd1 _12962_/A0 sky130_fd_sc_hd__buf_8
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1794 _17902_/Q vssd1 vssd1 vccd1 vccd1 _12756_/A sky130_fd_sc_hd__buf_12
X_19645_ _19645_/CLK _19645_/D vssd1 vssd1 vccd1 vccd1 _19645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16857_ _16836_/S _17923_/Q _16856_/X vssd1 vssd1 vccd1 vccd1 _17565_/B sky130_fd_sc_hd__o21ai_4
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15808_ _18600_/Q _15808_/A1 _15829_/S vssd1 vssd1 vccd1 vccd1 _18600_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16788_ _19284_/Q _16791_/C _16964_/A vssd1 vssd1 vccd1 vccd1 _16788_/Y sky130_fd_sc_hd__o21ai_1
X_19576_ _19608_/CLK _19576_/D vssd1 vssd1 vccd1 vccd1 _19576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18527_ _19286_/CLK _18527_/D vssd1 vssd1 vccd1 vccd1 _18527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15739_ _19484_/Q _15738_/X _15781_/S vssd1 vssd1 vccd1 vccd1 _15739_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ _10409_/A _09258_/X _09259_/X vssd1 vssd1 vccd1 vccd1 _09260_/X sky130_fd_sc_hd__a21o_1
XFILLER_244_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18458_ _19637_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09191_ _12442_/A _09643_/A vssd1 vssd1 vccd1 vccd1 _09191_/Y sky130_fd_sc_hd__nor2_1
X_17409_ _19493_/Q _17462_/B _17408_/X _17352_/A vssd1 vssd1 vccd1 vccd1 _19493_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18389_ _19465_/CLK _18389_/D vssd1 vssd1 vccd1 vccd1 _18389_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08975_ _08973_/X _08974_/X _11507_/S vssd1 vssd1 vccd1 vccd1 _08975_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09527_ _11172_/A1 _19560_/Q _09680_/B1 _19592_/Q vssd1 vssd1 vccd1 vccd1 _09527_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09458_ _10253_/A _10263_/A1 _19202_/Q _11406_/B2 vssd1 vssd1 vccd1 vccd1 _09458_/X
+ sky130_fd_sc_hd__a31o_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _18634_/Q _18056_/Q _09966_/S vssd1 vssd1 vccd1 vccd1 _09389_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11420_ _11498_/A1 _19208_/Q _19176_/Q _09290_/S vssd1 vssd1 vccd1 vccd1 _11420_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11351_ _11358_/A _11351_/B vssd1 vssd1 vccd1 vccd1 _11356_/A sky130_fd_sc_hd__and2_1
XFILLER_193_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10302_ _10747_/A1 _10301_/X _11501_/B1 vssd1 vssd1 vccd1 vccd1 _10302_/X sky130_fd_sc_hd__a21o_1
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14070_ _16488_/A0 _18012_/Q _14070_/S vssd1 vssd1 vccd1 vccd1 _18012_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ _11282_/A _11282_/B vssd1 vssd1 vccd1 vccd1 _11282_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13021_ _15872_/A _12506_/X _13010_/X _13020_/X _12510_/X vssd1 vssd1 vccd1 vccd1
+ _13023_/A sky130_fd_sc_hd__o221a_1
X_10233_ _10233_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__and2_2
XFILLER_3_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1002 _10414_/A2 vssd1 vssd1 vccd1 vccd1 _17685_/A0 sky130_fd_sc_hd__clkbuf_4
X_10164_ _17981_/Q _11447_/A2 _11371_/B1 vssd1 vssd1 vccd1 vccd1 _10164_/X sky130_fd_sc_hd__a21o_1
Xfanout1013 _15076_/S vssd1 vssd1 vccd1 vccd1 _15078_/S sky130_fd_sc_hd__buf_12
XFILLER_239_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1024 _16292_/A0 vssd1 vssd1 vccd1 vccd1 _16557_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1035 _15808_/A1 vssd1 vssd1 vccd1 vccd1 _16532_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 _08957_/Y vssd1 vssd1 vccd1 vccd1 _09523_/A sky130_fd_sc_hd__buf_12
X_10095_ _19065_/Q _19033_/Q _10168_/S vssd1 vssd1 vccd1 vccd1 _10095_/X sky130_fd_sc_hd__mux2_1
X_14972_ _17818_/Q _14982_/B vssd1 vssd1 vccd1 vccd1 _14972_/X sky130_fd_sc_hd__or2_1
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17760_ _19620_/CLK _17760_/D vssd1 vssd1 vccd1 vccd1 _17760_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1057 _15498_/S vssd1 vssd1 vccd1 vccd1 _15400_/S sky130_fd_sc_hd__buf_6
Xfanout1068 _12461_/Y vssd1 vssd1 vccd1 vccd1 _14033_/A1 sky130_fd_sc_hd__buf_4
XFILLER_266_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1079 _09995_/X vssd1 vssd1 vccd1 vccd1 _17659_/A0 sky130_fd_sc_hd__buf_6
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16711_ _19256_/Q _16717_/D _16710_/Y vssd1 vssd1 vccd1 vccd1 _19256_/D sky130_fd_sc_hd__o21a_1
XFILLER_208_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13923_ _19454_/Q _12582_/X _13922_/X vssd1 vssd1 vccd1 vccd1 _13923_/X sky130_fd_sc_hd__o21a_2
X_17691_ _17691_/A _17691_/B vssd1 vssd1 vccd1 vccd1 _17691_/Y sky130_fd_sc_hd__nand2_2
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16642_ _19236_/Q _16643_/C _16641_/Y vssd1 vssd1 vccd1 vccd1 _19236_/D sky130_fd_sc_hd__o21a_1
X_19430_ _19534_/CLK _19430_/D vssd1 vssd1 vccd1 vccd1 _19430_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13854_ _19324_/Q _13952_/A2 _13854_/B1 _13847_/X _13853_/X vssd1 vssd1 vccd1 vccd1
+ _13854_/Y sky130_fd_sc_hd__a2111oi_2
XFILLER_267_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12805_ _12668_/X _12673_/X _12821_/A vssd1 vssd1 vccd1 vccd1 _12805_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19361_ _19363_/CLK _19361_/D vssd1 vssd1 vccd1 vccd1 _19361_/Q sky130_fd_sc_hd__dfxtp_1
X_16573_ _16606_/A0 _19177_/Q _16585_/S vssd1 vssd1 vccd1 vccd1 _19177_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ _19386_/Q _13884_/A2 _13783_/X _13784_/X _13884_/C1 vssd1 vssd1 vccd1 vccd1
+ _13785_/X sky130_fd_sc_hd__o221a_4
X_10997_ _18550_/Q _11386_/S vssd1 vssd1 vccd1 vccd1 _10997_/X sky130_fd_sc_hd__or2_1
XFILLER_163_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18312_ _19608_/CLK _18312_/D vssd1 vssd1 vccd1 vccd1 _18312_/Q sky130_fd_sc_hd__dfxtp_1
X_15524_ _15516_/X _15517_/X _15523_/X _17540_/B1 _15633_/C1 vssd1 vssd1 vccd1 vccd1
+ _15524_/X sky130_fd_sc_hd__a221o_1
X_19292_ _19327_/CLK _19292_/D vssd1 vssd1 vccd1 vccd1 _19292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _12731_/X _12735_/Y _12933_/A vssd1 vssd1 vccd1 vccd1 _12988_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _19653_/A _18243_/D vssd1 vssd1 vccd1 vccd1 _18243_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15455_ _15455_/A _15455_/B vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__xnor2_2
X_12667_ _12756_/A _12740_/B vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__or2_4
XFILLER_129_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14406_ _17713_/A0 _18257_/Q _14416_/S vssd1 vssd1 vccd1 vccd1 _18257_/D sky130_fd_sc_hd__mux2_1
X_18174_ _19627_/CLK _18174_/D vssd1 vssd1 vccd1 vccd1 _18174_/Q sky130_fd_sc_hd__dfxtp_1
X_11618_ _11618_/A1 _18235_/Q _11613_/S _18970_/Q _11616_/S vssd1 vssd1 vccd1 vccd1
+ _11618_/X sky130_fd_sc_hd__o221a_1
X_15386_ _15387_/A _15387_/B vssd1 vssd1 vccd1 vccd1 _15386_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12598_ _12598_/A _12598_/B vssd1 vssd1 vccd1 vccd1 _12624_/A sky130_fd_sc_hd__or2_1
X_17125_ _19393_/Q _17120_/Y _17124_/X _14430_/B vssd1 vssd1 vccd1 vccd1 _19393_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14337_ _18194_/Q _16621_/A0 _14338_/S vssd1 vssd1 vccd1 vccd1 _18194_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11549_ _11550_/B _13797_/S _10380_/Y vssd1 vssd1 vccd1 vccd1 _11549_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17056_ _17123_/B _17074_/A2 _17055_/X _17378_/A vssd1 vssd1 vccd1 vccd1 _19361_/D
+ sky130_fd_sc_hd__o211a_1
X_14268_ _14268_/A _14268_/B vssd1 vssd1 vccd1 vccd1 _14268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16007_ _18719_/Q _16019_/A2 _16006_/X _14197_/A vssd1 vssd1 vccd1 vccd1 _18719_/D
+ sky130_fd_sc_hd__o211a_1
X_13219_ _13930_/A1 _13204_/X _13253_/B1 vssd1 vssd1 vccd1 vccd1 _13219_/X sky130_fd_sc_hd__o21a_1
X_14199_ _14203_/A _14199_/B vssd1 vssd1 vccd1 vccd1 _18097_/D sky130_fd_sc_hd__and2_1
XFILLER_140_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _17958_/CLK _17958_/D vssd1 vssd1 vccd1 vccd1 _17958_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_81_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19624_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_273_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1580 fanout1581/X vssd1 vssd1 vccd1 vccd1 _10356_/C1 sky130_fd_sc_hd__buf_6
X_16909_ _18758_/Q _16961_/A2 _16969_/B1 input222/X _16969_/C1 vssd1 vssd1 vccd1 vccd1
+ _16909_/X sky130_fd_sc_hd__a221o_2
Xfanout1591 _10211_/A1 vssd1 vssd1 vccd1 vccd1 _11503_/S1 sky130_fd_sc_hd__buf_6
XFILLER_39_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17889_ _17901_/CLK _17889_/D vssd1 vssd1 vccd1 vccd1 _17889_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19589_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19628_ _19628_/CLK _19628_/D vssd1 vssd1 vccd1 vccd1 _19628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19559_ _19591_/CLK _19559_/D vssd1 vssd1 vccd1 vccd1 _19559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09312_ _11417_/B1 _09310_/X _09311_/X _09297_/X vssd1 vssd1 vccd1 vccd1 _09312_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09243_ _09652_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09243_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09174_ _11017_/A1 _19628_/Q _18917_/Q _09344_/S vssd1 vssd1 vccd1 vccd1 _09174_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput105 dout0[8] vssd1 vssd1 vccd1 vccd1 input105/X sky130_fd_sc_hd__clkbuf_2
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput116 dout1[18] vssd1 vssd1 vccd1 vccd1 input116/X sky130_fd_sc_hd__clkbuf_2
XFILLER_276_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput127 dout1[28] vssd1 vssd1 vccd1 vccd1 input127/X sky130_fd_sc_hd__clkbuf_2
XFILLER_276_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput138 dout1[38] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_hd__buf_2
X_08958_ _08958_/A _08958_/B vssd1 vssd1 vccd1 vccd1 _08958_/X sky130_fd_sc_hd__or2_4
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput149 dout1[48] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_hd__buf_2
XFILLER_236_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ _12267_/A _17891_/Q _17890_/Q vssd1 vssd1 vccd1 vccd1 _12439_/A sky130_fd_sc_hd__or3b_4
XFILLER_57_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ _10785_/A _10918_/X _10919_/X _11570_/B1 vssd1 vssd1 vccd1 vccd1 _10920_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10851_ _10785_/A _10849_/X _10850_/X _11563_/B1 vssd1 vssd1 vccd1 vccd1 _10851_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_271_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ _11673_/B _13912_/B1 _13912_/A2 _10984_/A _14153_/A vssd1 vssd1 vccd1 vccd1
+ _13570_/X sky130_fd_sc_hd__a221o_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10782_ _11305_/A1 _18225_/Q _11302_/S _18960_/Q vssd1 vssd1 vccd1 vccd1 _10782_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_198_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12521_ _19522_/Q _12771_/A _12580_/A vssd1 vssd1 vccd1 vccd1 _12521_/X sky130_fd_sc_hd__and3_1
XFILLER_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _14220_/A _15786_/A2 _15239_/Y _12318_/A vssd1 vssd1 vccd1 vccd1 _15243_/A
+ sky130_fd_sc_hd__o22a_4
X_12452_ _12755_/A _12587_/B vssd1 vssd1 vccd1 vccd1 _12452_/Y sky130_fd_sc_hd__nand2_1
X_11403_ _18856_/Q _18888_/Q _11403_/S vssd1 vssd1 vccd1 vccd1 _11403_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15171_ _15171_/A _15171_/B vssd1 vssd1 vccd1 vccd1 _15179_/A sky130_fd_sc_hd__nand2_1
X_12383_ _17902_/Q _12382_/A _12382_/Y _12383_/C1 vssd1 vssd1 vccd1 vccd1 _17902_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14122_ _16539_/A0 _18061_/Q _14139_/S vssd1 vssd1 vccd1 vccd1 _18061_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11334_ _11488_/A _11828_/A vssd1 vssd1 vccd1 vccd1 _11334_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14053_ _17703_/A0 _17995_/Q _14072_/S vssd1 vssd1 vccd1 vccd1 _17995_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18930_ _19641_/CLK _18930_/D vssd1 vssd1 vccd1 vccd1 _18930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ _11263_/X _11264_/X _11285_/S vssd1 vssd1 vccd1 vccd1 _11265_/X sky130_fd_sc_hd__mux2_1
XFILLER_268_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13004_ _12987_/Y _13003_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _13004_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_279_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10216_ _10214_/X _10215_/X _10225_/S vssd1 vssd1 vccd1 vccd1 _10216_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18861_ _19075_/CLK _18861_/D vssd1 vssd1 vccd1 vccd1 _18861_/Q sky130_fd_sc_hd__dfxtp_1
X_11196_ _11277_/A1 _19211_/Q _19179_/Q _10717_/S vssd1 vssd1 vccd1 vccd1 _11196_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_267_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17812_ _19492_/CLK _17812_/D vssd1 vssd1 vccd1 vccd1 _17812_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _09708_/A _10142_/X _10146_/X _08895_/A vssd1 vssd1 vccd1 vccd1 _10147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18792_ _19208_/CLK _18792_/D vssd1 vssd1 vccd1 vccd1 _18792_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14955_ _18127_/Q _14994_/B _14934_/X _14954_/X vssd1 vssd1 vccd1 vccd1 _14955_/X
+ sky130_fd_sc_hd__o211a_1
X_17743_ _18643_/Q vssd1 vssd1 vccd1 vccd1 _18643_/D sky130_fd_sc_hd__clkbuf_2
X_10078_ _11750_/A _11750_/B _13195_/S vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__a21boi_4
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13906_ _17949_/Q _13973_/A2 _13904_/Y _13905_/X _14342_/A vssd1 vssd1 vccd1 vccd1
+ _17949_/D sky130_fd_sc_hd__o221a_1
XFILLER_208_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14886_ input53/X input89/X _14947_/S vssd1 vssd1 vccd1 vccd1 _14887_/A sky130_fd_sc_hd__mux2_2
X_17674_ _17674_/A0 _19601_/Q _17690_/S vssd1 vssd1 vccd1 vccd1 _19601_/D sky130_fd_sc_hd__mux2_1
XFILLER_263_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19413_ _19477_/CLK _19413_/D vssd1 vssd1 vccd1 vccd1 _19413_/Q sky130_fd_sc_hd__dfxtp_2
X_16625_ _19228_/Q input248/X _16627_/S vssd1 vssd1 vccd1 vccd1 _19228_/D sky130_fd_sc_hd__mux2_1
X_13837_ _18128_/Q _13837_/B vssd1 vssd1 vccd1 vccd1 _13838_/B sky130_fd_sc_hd__nor2_1
XFILLER_262_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16556_ _16622_/A0 _19161_/Q _16556_/S vssd1 vssd1 vccd1 vccd1 _19161_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19344_ _19543_/CLK _19344_/D vssd1 vssd1 vccd1 vccd1 _19344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13768_ _13761_/X _13764_/Y _13766_/X _13767_/X vssd1 vssd1 vccd1 vccd1 _13768_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12719_ _13314_/S _12719_/B vssd1 vssd1 vccd1 vccd1 _12719_/X sky130_fd_sc_hd__or2_1
X_15507_ _15554_/A vssd1 vssd1 vccd1 vccd1 _15511_/A sky130_fd_sc_hd__inv_2
X_19275_ _19276_/CLK _19275_/D vssd1 vssd1 vccd1 vccd1 _19275_/Q sky130_fd_sc_hd__dfxtp_1
X_16487_ _16553_/A0 _19094_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _19094_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13699_ _11541_/A _13912_/A2 _12836_/Y _13697_/A _14153_/A vssd1 vssd1 vccd1 vccd1
+ _13699_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15438_ _19439_/Q _15124_/B _17166_/A vssd1 vssd1 vccd1 vccd1 _15438_/Y sky130_fd_sc_hd__o21ai_1
X_18226_ _19602_/CLK _18226_/D vssd1 vssd1 vccd1 vccd1 _18226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18157_ _19642_/CLK _18157_/D vssd1 vssd1 vccd1 vccd1 _18157_/Q sky130_fd_sc_hd__dfxtp_1
X_15369_ _15369_/A _15385_/B _15369_/C vssd1 vssd1 vccd1 vccd1 _15369_/X sky130_fd_sc_hd__and3_1
XFILLER_190_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17108_ _17202_/B _17108_/A2 _17107_/X _17366_/A vssd1 vssd1 vccd1 vccd1 _19387_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18088_ _18749_/CLK _18088_/D vssd1 vssd1 vccd1 vccd1 _18088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09930_ _10262_/A1 _18134_/Q _18780_/Q _11472_/C _11397_/A1 vssd1 vssd1 vccd1 vccd1
+ _09930_/X sky130_fd_sc_hd__a221o_1
X_17039_ _19356_/Q _17041_/B vssd1 vssd1 vccd1 vccd1 _17039_/X sky130_fd_sc_hd__or2_1
XFILLER_113_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout806 _15817_/S vssd1 vssd1 vccd1 vccd1 _15829_/S sky130_fd_sc_hd__buf_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _17897_/Q _15120_/A vssd1 vssd1 vccd1 vccd1 _09861_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout817 _14325_/S vssd1 vssd1 vccd1 vccd1 _14339_/S sky130_fd_sc_hd__buf_12
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout828 _12019_/S vssd1 vssd1 vccd1 vccd1 _12021_/S sky130_fd_sc_hd__buf_12
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout839 _17710_/A0 vssd1 vssd1 vccd1 vccd1 _17644_/A0 sky130_fd_sc_hd__clkbuf_2
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _18442_/Q _18343_/Q _09797_/S vssd1 vssd1 vccd1 vccd1 _09792_/X sky130_fd_sc_hd__mux2_1
XFILLER_218_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09226_ _09946_/B1 _15303_/A _09193_/X vssd1 vssd1 vccd1 vccd1 _12599_/B sky130_fd_sc_hd__o21a_4
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09157_ _09049_/Y _09156_/X _09152_/X _09030_/X vssd1 vssd1 vccd1 vccd1 _09157_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_257_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _12408_/A _09285_/C vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__and2_4
XFILLER_174_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11050_ _11428_/A _11049_/X _11417_/B1 vssd1 vssd1 vccd1 vccd1 _11050_/X sky130_fd_sc_hd__a21o_1
XFILLER_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10001_ _18626_/Q _18048_/Q _10001_/S vssd1 vssd1 vccd1 vccd1 _10001_/X sky130_fd_sc_hd__mux2_1
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _18475_/Q _14889_/B1 _14739_/Y _17330_/A vssd1 vssd1 vccd1 vccd1 _18475_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _11666_/A _11952_/A2 _11774_/B _11663_/A vssd1 vssd1 vccd1 vccd1 _14342_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903_ _11365_/B2 _14510_/A0 _10902_/X _11133_/B2 vssd1 vssd1 vccd1 vccd1 _13581_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_260_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _14671_/A _14680_/C vssd1 vssd1 vccd1 vccd1 _14671_/X sky130_fd_sc_hd__or2_2
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11883_ _10415_/B _11864_/B _11887_/B1 vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__o21ai_2
XFILLER_264_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _16608_/A0 _19019_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _19019_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13622_ _13622_/A _13622_/B vssd1 vssd1 vccd1 vccd1 _13622_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10834_ _11141_/A _10834_/B vssd1 vssd1 vccd1 vccd1 _10834_/Y sky130_fd_sc_hd__nor2_1
X_17390_ _17523_/B vssd1 vssd1 vccd1 vccd1 _17390_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_260_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16341_ _18953_/Q _16540_/A0 _16358_/S vssd1 vssd1 vccd1 vccd1 _18953_/D sky130_fd_sc_hd__mux2_1
X_13553_ _19541_/Q _13946_/B vssd1 vssd1 vccd1 vccd1 _13553_/X sky130_fd_sc_hd__or2_1
XFILLER_213_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10765_ _19056_/Q _19024_/Q _10864_/S vssd1 vssd1 vccd1 vccd1 _10765_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12504_ _12572_/A _12572_/B _12572_/C _12503_/Y vssd1 vssd1 vccd1 vccd1 _13165_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_157_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19060_ _19609_/CLK _19060_/D vssd1 vssd1 vccd1 vccd1 _19060_/Q sky130_fd_sc_hd__dfxtp_1
X_16272_ _09105_/A _18886_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _18886_/D sky130_fd_sc_hd__mux2_1
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ _11214_/A _11212_/Y _13466_/A vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__o21bai_1
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10696_ _11480_/C1 _10693_/X _10695_/X vssd1 vssd1 vccd1 vccd1 _10696_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18011_ _19613_/CLK _18011_/D vssd1 vssd1 vccd1 vccd1 _18011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15223_ _15223_/A _15223_/B vssd1 vssd1 vccd1 vccd1 _15236_/B sky130_fd_sc_hd__nor2_1
XFILLER_201_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12435_ _12435_/A _13260_/A vssd1 vssd1 vccd1 vccd1 _12587_/B sky130_fd_sc_hd__nor2_8
XFILLER_218_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15154_ _15155_/A _15155_/B vssd1 vssd1 vccd1 vccd1 _15171_/A sky130_fd_sc_hd__or2_2
X_12366_ _18382_/Q _12417_/B1 _09243_/Y _08858_/A vssd1 vssd1 vccd1 vccd1 _12367_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput409 _18503_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_ack_o sky130_fd_sc_hd__buf_4
XFILLER_126_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14105_ _17688_/A0 _18045_/Q _14106_/S vssd1 vssd1 vccd1 vccd1 _18045_/D sky130_fd_sc_hd__mux2_1
XFILLER_271_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11317_ _19049_/Q _19017_/Q _11325_/S vssd1 vssd1 vccd1 vccd1 _11317_/X sky130_fd_sc_hd__mux2_1
X_15085_ _19383_/Q _15092_/B _15085_/C vssd1 vssd1 vccd1 vccd1 _15085_/X sky130_fd_sc_hd__and3_1
XFILLER_181_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12297_ _18084_/Q _12277_/B _14692_/A2 _18507_/Q vssd1 vssd1 vccd1 vccd1 _14675_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18913_ _19624_/CLK _18913_/D vssd1 vssd1 vccd1 vccd1 _18913_/Q sky130_fd_sc_hd__dfxtp_1
X_14036_ _14036_/A _14036_/B vssd1 vssd1 vccd1 vccd1 _14036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11248_ _11246_/X _11247_/X _11248_/S vssd1 vssd1 vccd1 vccd1 _11248_/X sky130_fd_sc_hd__mux2_1
XFILLER_268_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18844_ _19201_/CLK _18844_/D vssd1 vssd1 vccd1 vccd1 _18844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11179_ _11332_/B1 _11177_/X _11178_/X vssd1 vssd1 vccd1 vccd1 _11837_/A sky130_fd_sc_hd__o21ai_4
XFILLER_255_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18775_ _18775_/CLK _18775_/D vssd1 vssd1 vccd1 vccd1 _18775_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _18709_/Q _16005_/A2 _15986_/X _14197_/A vssd1 vssd1 vccd1 vccd1 _18709_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_208_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17726_ _18626_/Q vssd1 vssd1 vccd1 vccd1 _18626_/D sky130_fd_sc_hd__clkbuf_2
X_14938_ _14938_/A vssd1 vssd1 vccd1 vccd1 _14938_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17657_ _17690_/A0 _19585_/Q _17657_/S vssd1 vssd1 vccd1 vccd1 _19585_/D sky130_fd_sc_hd__mux2_1
XFILLER_224_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14869_ _14865_/Y _14868_/X _14879_/B1 vssd1 vssd1 vccd1 vccd1 _14869_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_24_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16608_ _16608_/A0 _19211_/Q _16619_/S vssd1 vssd1 vccd1 vccd1 _19211_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17588_ _19536_/Q _17561_/B _17588_/B1 _17587_/X vssd1 vssd1 vccd1 vccd1 _19536_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_251_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19327_ _19327_/CLK _19327_/D vssd1 vssd1 vccd1 vccd1 _19327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16539_ _16539_/A0 _19144_/Q _16556_/S vssd1 vssd1 vccd1 vccd1 _19144_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19258_ _19261_/CLK _19258_/D vssd1 vssd1 vccd1 vccd1 _19258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09011_ input168/X input139/X _09990_/S vssd1 vssd1 vccd1 vccd1 _09012_/C sky130_fd_sc_hd__mux2_8
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18209_ _19591_/CLK _18209_/D vssd1 vssd1 vccd1 vccd1 _18209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19189_ _19644_/CLK _19189_/D vssd1 vssd1 vccd1 vccd1 _19189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09913_ _09457_/B _18017_/Q _17985_/Q _11167_/B _10337_/S1 vssd1 vssd1 vccd1 vccd1
+ _09913_/X sky130_fd_sc_hd__o221a_1
Xfanout603 _17475_/A2 vssd1 vssd1 vccd1 vccd1 _17520_/A2 sky130_fd_sc_hd__buf_4
Xfanout614 _17622_/A2 vssd1 vssd1 vccd1 vccd1 _17624_/A2 sky130_fd_sc_hd__buf_4
XFILLER_101_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout625 _16980_/X vssd1 vssd1 vccd1 vccd1 _17008_/A2 sky130_fd_sc_hd__buf_4
Xfanout636 _17589_/B vssd1 vssd1 vccd1 vccd1 _17583_/B sky130_fd_sc_hd__buf_4
X_09844_ _19101_/Q _19133_/Q _11147_/S vssd1 vssd1 vccd1 vccd1 _09844_/X sky130_fd_sc_hd__mux2_1
Xfanout647 _17073_/B vssd1 vssd1 vccd1 vccd1 _17107_/B sky130_fd_sc_hd__buf_4
XFILLER_258_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout658 _13781_/B1 vssd1 vssd1 vccd1 vccd1 _13947_/B1 sky130_fd_sc_hd__buf_4
XFILLER_274_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout669 _11846_/A vssd1 vssd1 vccd1 vccd1 _11859_/A sky130_fd_sc_hd__buf_12
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09775_ _11790_/B _11790_/C _11790_/D _15120_/A vssd1 vssd1 vccd1 vccd1 _09775_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_274_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ _11312_/A1 _19578_/Q _09108_/B _19610_/Q vssd1 vssd1 vccd1 vccd1 _10550_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_183_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _10747_/A1 _09208_/X _09204_/X _11501_/B1 vssd1 vssd1 vccd1 vccd1 _09209_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_167_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10481_ _11566_/A1 _19156_/Q _10840_/S _19124_/Q vssd1 vssd1 vccd1 vccd1 _10481_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_120_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12220_ _17871_/Q _12218_/B _12219_/Y vssd1 vssd1 vccd1 vccd1 _17871_/D sky130_fd_sc_hd__o21a_1
XFILLER_182_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12151_ _17845_/Q _12152_/C _17846_/Q vssd1 vssd1 vccd1 vccd1 _12153_/B sky130_fd_sc_hd__a21oi_1
XFILLER_163_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11102_ _11332_/B1 _11100_/X _11101_/X vssd1 vssd1 vccd1 vccd1 _11841_/A sky130_fd_sc_hd__o21ai_2
XFILLER_123_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ _17916_/Q _12088_/A2 _12081_/X _17328_/A vssd1 vssd1 vccd1 vccd1 _17818_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15910_ _18679_/Q _15910_/A2 _15909_/X _15910_/C1 vssd1 vssd1 vccd1 vccd1 _18679_/D
+ sky130_fd_sc_hd__o211a_1
X_11033_ _18644_/Q _18066_/Q _19085_/Q _18989_/Q _11426_/B2 _11510_/S1 vssd1 vssd1
+ vccd1 vccd1 _11034_/B sky130_fd_sc_hd__mux4_1
XFILLER_2_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16890_ _16970_/A1 _17931_/Q _16889_/X vssd1 vssd1 vccd1 vccd1 _17581_/A sky130_fd_sc_hd__o21a_4
XFILLER_1_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _18659_/Q _15843_/A _15840_/Y _14177_/A vssd1 vssd1 vccd1 vccd1 _18659_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_209_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18660_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_253_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _19159_/CLK _18560_/D vssd1 vssd1 vccd1 vccd1 _18560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _18592_/Q _15772_/B vssd1 vssd1 vccd1 vccd1 _15772_/X sky130_fd_sc_hd__or2_1
X_12984_ _13462_/A _12979_/X _12980_/Y _12983_/X vssd1 vssd1 vccd1 vccd1 _12984_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_264_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _18586_/Q _17527_/A1 _17516_/C1 vssd1 vssd1 vccd1 vccd1 _17511_/X sky130_fd_sc_hd__o21a_1
XFILLER_245_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14723_ _17793_/Q _14722_/X _14993_/S vssd1 vssd1 vccd1 vccd1 _14723_/X sky130_fd_sc_hd__mux2_1
X_11935_ _11959_/B2 _11836_/B _11935_/B1 input221/X vssd1 vssd1 vccd1 vccd1 _11935_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_245_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18491_ _19285_/CLK _18491_/D vssd1 vssd1 vccd1 vccd1 _18491_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_530 _11853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_541 _18113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14654_ _17713_/A0 _18460_/Q _14664_/S vssd1 vssd1 vccd1 vccd1 _18460_/D sky130_fd_sc_hd__mux2_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _18111_/Q _17463_/A2 _17440_/X _17441_/X vssd1 vssd1 vccd1 vccd1 _17442_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11866_ _14141_/B _11828_/X _11865_/Y _11859_/B vssd1 vssd1 vccd1 vccd1 _11866_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13323_/B _13603_/X _13604_/X _13323_/X vssd1 vssd1 vccd1 vccd1 _13605_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10817_ _10817_/A1 _18154_/Q _18800_/Q _11360_/B2 vssd1 vssd1 vccd1 vccd1 _10817_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14585_ _18401_/Q _14589_/A2 _14589_/B1 input30/X vssd1 vssd1 vccd1 vccd1 _14586_/B
+ sky130_fd_sc_hd__o22a_1
X_17373_ _19484_/Q _17205_/B _17379_/S vssd1 vssd1 vccd1 vccd1 _17374_/B sky130_fd_sc_hd__mux2_1
X_11797_ _11799_/A _11799_/B _11825_/B vssd1 vssd1 vccd1 vccd1 _11797_/X sky130_fd_sc_hd__and3_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19112_ _19630_/CLK _19112_/D vssd1 vssd1 vccd1 vccd1 _19112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16324_ _17722_/A0 _18937_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _18937_/D sky130_fd_sc_hd__mux2_1
X_13536_ _13962_/B _13535_/X _11062_/B vssd1 vssd1 vccd1 vccd1 _13536_/X sky130_fd_sc_hd__a21o_1
X_10748_ _10741_/X _10747_/X _10731_/X vssd1 vssd1 vccd1 vccd1 _10748_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19043_ _19594_/CLK _19043_/D vssd1 vssd1 vccd1 vccd1 _19043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16255_ _17719_/A0 _18870_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _18870_/D sky130_fd_sc_hd__mux2_1
X_13467_ _13486_/A1 _14145_/B _13909_/B1 vssd1 vssd1 vccd1 vccd1 _13467_/Y sky130_fd_sc_hd__a21oi_1
X_10679_ _11556_/C _10679_/B vssd1 vssd1 vccd1 vccd1 _10679_/Y sky130_fd_sc_hd__nor2_2
XFILLER_127_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _18567_/Q _15224_/C vssd1 vssd1 vccd1 vccd1 _15206_/X sky130_fd_sc_hd__xor2_1
X_12418_ _12427_/A _12418_/B vssd1 vssd1 vccd1 vccd1 _12418_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16186_ _16418_/A0 _18803_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _18803_/D sky130_fd_sc_hd__mux2_1
X_13398_ _18114_/Q _13397_/C _18115_/Q vssd1 vssd1 vccd1 vccd1 _13399_/B sky130_fd_sc_hd__a21oi_1
XFILLER_182_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15137_ _15137_/A _15137_/B vssd1 vssd1 vccd1 vccd1 _15138_/C sky130_fd_sc_hd__and2_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12349_ _12349_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _12349_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15068_ _18552_/Q _16314_/A0 _15079_/S vssd1 vssd1 vccd1 vccd1 _18552_/D sky130_fd_sc_hd__mux2_1
X_14019_ _14033_/A1 _13659_/X _14018_/X _14417_/A vssd1 vssd1 vccd1 vccd1 _17974_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18827_ _19634_/CLK _18827_/D vssd1 vssd1 vccd1 vccd1 _18827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09560_ _12613_/B _09561_/B vssd1 vssd1 vccd1 vccd1 _09560_/X sky130_fd_sc_hd__and2_2
X_18758_ _18761_/CLK _18758_/D vssd1 vssd1 vccd1 vccd1 _18758_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_237_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17709_ _17709_/A0 _19635_/Q _17723_/S vssd1 vssd1 vccd1 vccd1 _19635_/D sky130_fd_sc_hd__mux2_1
XFILLER_247_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09491_ _17958_/Q _11216_/A2 _08947_/X _17926_/Q _09490_/X vssd1 vssd1 vccd1 vccd1
+ _09491_/X sky130_fd_sc_hd__a221o_2
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18689_ _18691_/CLK _18689_/D vssd1 vssd1 vccd1 vccd1 _18689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1409 fanout1415/X vssd1 vssd1 vccd1 vccd1 _10168_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_274_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09827_ _18441_/Q _10001_/S _10004_/A1 _09826_/X vssd1 vssd1 vccd1 vccd1 _09827_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_246_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout488 _14950_/B1 vssd1 vssd1 vccd1 vccd1 _14879_/B1 sky130_fd_sc_hd__buf_12
XFILLER_150_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout499 _11919_/X vssd1 vssd1 vccd1 vccd1 _11949_/B1 sky130_fd_sc_hd__buf_4
XFILLER_86_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09758_ _09756_/X _09757_/X _11562_/S vssd1 vssd1 vccd1 vccd1 _09758_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _09687_/X _09688_/X _11161_/S vssd1 vssd1 vccd1 vccd1 _09690_/B sky130_fd_sc_hd__mux2_1
XFILLER_15_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11968_/B2 _11919_/B vssd1 vssd1 vccd1 vccd1 _11720_/X sky130_fd_sc_hd__and2b_4
XFILLER_14_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11651_ _14141_/A _11651_/B vssd1 vssd1 vccd1 vccd1 _11653_/B sky130_fd_sc_hd__nor2_1
XFILLER_230_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10602_ _10602_/A _12650_/B vssd1 vssd1 vccd1 vccd1 _10603_/B sky130_fd_sc_hd__nor2_4
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14370_ _18222_/Q _17644_/A0 _14380_/S vssd1 vssd1 vccd1 vccd1 _18222_/D sky130_fd_sc_hd__mux2_1
X_11582_ _10471_/S _11581_/X _11580_/X vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__o21ai_1
XFILLER_196_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ _13931_/A _13321_/B _13321_/C vssd1 vssd1 vccd1 vccd1 _13321_/X sky130_fd_sc_hd__or3_1
X_10533_ _18463_/Q _18364_/Q _10613_/S vssd1 vssd1 vccd1 vccd1 _10533_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ _18741_/Q _18740_/Q vssd1 vssd1 vccd1 vccd1 _16063_/B sky130_fd_sc_hd__nand2_2
XFILLER_182_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13252_ _12455_/Y _13251_/X _13238_/X vssd1 vssd1 vccd1 vccd1 _13252_/X sky130_fd_sc_hd__a21o_1
X_10464_ _10625_/A1 _19220_/Q _19188_/Q _10613_/S _09095_/A vssd1 vssd1 vccd1 vccd1
+ _10464_/X sky130_fd_sc_hd__a221o_1
XFILLER_89_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ _12203_/A _12208_/C vssd1 vssd1 vccd1 vccd1 _12203_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _12586_/X _13163_/Y _13563_/B1 vssd1 vssd1 vccd1 vccd1 _13183_/X sky130_fd_sc_hd__a21o_1
X_10395_ _18869_/Q _18901_/Q _10864_/S vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__mux2_1
X_12134_ _17839_/Q _12136_/C _12133_/Y vssd1 vssd1 vccd1 vccd1 _17839_/D sky130_fd_sc_hd__o21a_1
XFILLER_269_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17991_ _18880_/CLK _17991_/D vssd1 vssd1 vccd1 vccd1 _17991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16942_ _16848_/S _17944_/Q _16941_/X vssd1 vssd1 vccd1 vccd1 _17193_/B sky130_fd_sc_hd__o21a_4
Xfanout1910 input205/X vssd1 vssd1 vccd1 vccd1 _11712_/A sky130_fd_sc_hd__buf_4
X_12065_ _17810_/Q _12085_/B vssd1 vssd1 vccd1 vccd1 _12065_/X sky130_fd_sc_hd__or2_1
XFILLER_123_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11016_ _18861_/Q _18893_/Q _11395_/C vssd1 vssd1 vccd1 vccd1 _11016_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16873_ _18749_/Q _12276_/A _16877_/B1 input244/X _12483_/A vssd1 vssd1 vccd1 vccd1
+ _16873_/X sky130_fd_sc_hd__a221o_1
XFILLER_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18612_ _19636_/CLK _18612_/D vssd1 vssd1 vccd1 vccd1 _18612_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15824_ _18616_/Q _17714_/A0 _15829_/S vssd1 vssd1 vccd1 vccd1 _18616_/D sky130_fd_sc_hd__mux2_1
XFILLER_219_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ _19592_/CLK _19592_/D vssd1 vssd1 vccd1 vccd1 _19592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _18543_/CLK _18543_/D vssd1 vssd1 vccd1 vccd1 _18543_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12967_ _19300_/Q _13952_/A2 _12551_/Y vssd1 vssd1 vccd1 vccd1 _12967_/X sky130_fd_sc_hd__a21o_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15755_ _15753_/Y _15755_/B vssd1 vssd1 vccd1 vccd1 _15758_/A sky130_fd_sc_hd__nand2b_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14706_ _18659_/Q _16819_/B _14685_/X _14875_/A1 _14705_/X vssd1 vssd1 vccd1 vccd1
+ _14706_/X sky130_fd_sc_hd__a311o_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _18572_/Q _11918_/A2 _11664_/X _13224_/A vssd1 vssd1 vccd1 vccd1 _11918_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_261_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18474_ _19464_/CLK _18474_/D vssd1 vssd1 vccd1 vccd1 _18474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_261_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_360 _11252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15686_ _15686_/A _15686_/B vssd1 vssd1 vccd1 vccd1 _15686_/X sky130_fd_sc_hd__or2_1
X_12898_ _13896_/B2 _12891_/X _12897_/X _12732_/S vssd1 vssd1 vccd1 vccd1 _12898_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_371 _18274_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_382 _15854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17425_ _13125_/A _17445_/A2 _15117_/A _17797_/Q _17445_/C1 vssd1 vssd1 vccd1 vccd1
+ _17425_/X sky130_fd_sc_hd__a221o_1
XFILLER_178_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_393 _09004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14637_ _17696_/A0 _18443_/Q _14660_/S vssd1 vssd1 vccd1 vccd1 _18443_/D sky130_fd_sc_hd__mux2_1
X_11849_ _11909_/A _11849_/B vssd1 vssd1 vccd1 vccd1 _11849_/X sky130_fd_sc_hd__and2_1
XFILLER_221_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17356_ _17356_/A _17356_/B vssd1 vssd1 vccd1 vccd1 _19475_/D sky130_fd_sc_hd__and2_1
X_14568_ _14576_/A _14568_/B vssd1 vssd1 vccd1 vccd1 _18392_/D sky130_fd_sc_hd__or2_1
XFILLER_158_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19619_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16307_ _17705_/A0 _18920_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _18920_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13519_ _17873_/Q _13747_/A2 _13518_/X _13747_/B2 vssd1 vssd1 vccd1 vccd1 _13519_/X
+ sky130_fd_sc_hd__a22o_1
X_14499_ _17701_/A0 _18349_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _18349_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17287_ _18123_/Q _15717_/B2 _17503_/A _17313_/B vssd1 vssd1 vccd1 vccd1 _17287_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_256_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19026_ _19219_/CLK _19026_/D vssd1 vssd1 vccd1 vccd1 _19026_/Q sky130_fd_sc_hd__dfxtp_1
X_16238_ _16602_/A0 _18853_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _18853_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16169_ _17666_/A0 _18786_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _18786_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08991_ _08991_/A _17796_/Q _17794_/Q _17795_/Q vssd1 vssd1 vccd1 vccd1 _08991_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_142_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09612_ _18537_/Q _18412_/Q _18021_/Q _17989_/Q _10313_/S _10266_/S1 vssd1 vssd1
+ vccd1 vccd1 _09612_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09543_ _09541_/X _09542_/X _09845_/S vssd1 vssd1 vccd1 vccd1 _09544_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09474_ _12612_/B _09475_/B vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__and2_4
XFILLER_240_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10180_ _10180_/A _10180_/B vssd1 vssd1 vccd1 vccd1 _10180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1206 _12753_/X vssd1 vssd1 vccd1 vccd1 _14156_/A0 sky130_fd_sc_hd__buf_6
XFILLER_266_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1217 _12442_/D vssd1 vssd1 vccd1 vccd1 _13602_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1228 _12318_/A vssd1 vssd1 vccd1 vccd1 _15481_/B sky130_fd_sc_hd__buf_2
XFILLER_278_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1239 _11257_/C1 vssd1 vssd1 vccd1 vccd1 _11800_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_275_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ _13904_/A _13870_/B vssd1 vssd1 vccd1 vccd1 _13870_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12821_ _12821_/A _12821_/B vssd1 vssd1 vccd1 vccd1 _12821_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ _19475_/Q _19409_/Q vssd1 vssd1 vccd1 vccd1 _15540_/Y sky130_fd_sc_hd__nor2_1
X_12752_ _13315_/S _12751_/Y _13197_/B1 vssd1 vssd1 vccd1 vccd1 _12752_/X sky130_fd_sc_hd__a21o_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11703_ _11706_/C _11706_/B _11702_/X _18268_/Q vssd1 vssd1 vccd1 vccd1 _14345_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _19472_/Q _19406_/Q vssd1 vssd1 vccd1 vccd1 _15472_/B sky130_fd_sc_hd__or2_1
X_12683_ _12942_/S _12872_/B vssd1 vssd1 vccd1 vccd1 _12683_/X sky130_fd_sc_hd__or2_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17210_/A _17210_/B vssd1 vssd1 vccd1 vccd1 _19421_/D sky130_fd_sc_hd__nor2_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _11721_/Y _18274_/D vssd1 vssd1 vccd1 vccd1 _18273_/D sky130_fd_sc_hd__and2b_1
X_11634_ _11634_/A _11634_/B vssd1 vssd1 vccd1 vccd1 _13891_/A sky130_fd_sc_hd__or2_4
X_18190_ _19643_/CLK _18190_/D vssd1 vssd1 vccd1 vccd1 _18190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14353_ _18205_/Q _16461_/A0 _14380_/S vssd1 vssd1 vccd1 vccd1 _18205_/D sky130_fd_sc_hd__mux2_1
X_17141_ _17141_/A _17141_/B vssd1 vssd1 vccd1 vccd1 _19398_/D sky130_fd_sc_hd__nor2_1
X_11565_ _11565_/A1 _18235_/Q _11070_/S _18970_/Q vssd1 vssd1 vccd1 vccd1 _11565_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _19308_/Q _12583_/Y _13302_/X _13303_/X vssd1 vssd1 vccd1 vccd1 _13304_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_196_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10516_ _19643_/Q _18932_/Q _10582_/S vssd1 vssd1 vccd1 vccd1 _10516_/X sky130_fd_sc_hd__mux2_1
X_17072_ _17577_/A _17108_/A2 _17071_/X _17469_/C1 vssd1 vssd1 vccd1 vccd1 _19369_/D
+ sky130_fd_sc_hd__o211a_1
X_14284_ _16602_/A0 _18143_/Q _14304_/S vssd1 vssd1 vccd1 vccd1 _18143_/D sky130_fd_sc_hd__mux2_1
X_11496_ _10419_/S _11491_/X _11495_/X vssd1 vssd1 vccd1 vccd1 _11496_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16023_ _16020_/Y _16022_/X _16021_/X _16052_/A vssd1 vssd1 vccd1 vccd1 _18726_/D
+ sky130_fd_sc_hd__o211a_1
X_13235_ _18111_/Q _13271_/C vssd1 vssd1 vccd1 vccd1 _13236_/A sky130_fd_sc_hd__xnor2_2
X_10447_ _11602_/C1 _10440_/X _11286_/B1 vssd1 vssd1 vccd1 vccd1 _10447_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_237_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13166_ _19240_/Q _13425_/A2 _13425_/B1 _19272_/Q vssd1 vssd1 vccd1 vccd1 _13166_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10378_ _18128_/Q _10377_/Y _13739_/A vssd1 vssd1 vccd1 vccd1 _12653_/B sky130_fd_sc_hd__mux2_8
XFILLER_151_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12117_ _17833_/Q _12120_/C _16811_/A vssd1 vssd1 vccd1 vccd1 _12117_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_153_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19399_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_269_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17974_ _17975_/CLK _17974_/D vssd1 vssd1 vccd1 vccd1 _17974_/Q sky130_fd_sc_hd__dfxtp_1
X_13097_ _11742_/B _13912_/B1 _13096_/X vssd1 vssd1 vccd1 vccd1 _13097_/X sky130_fd_sc_hd__a21bo_1
X_16925_ _18762_/Q _16965_/A2 _16965_/B1 input227/X _16965_/C1 vssd1 vssd1 vccd1 vccd1
+ _16925_/X sky130_fd_sc_hd__a221o_2
Xfanout1740 _18274_/Q vssd1 vssd1 vccd1 vccd1 _15009_/A1 sky130_fd_sc_hd__clkbuf_4
X_12048_ _17899_/Q _12052_/A2 _12047_/X _13100_/A vssd1 vssd1 vccd1 vccd1 _17801_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1751 _17919_/Q vssd1 vssd1 vccd1 vccd1 _15549_/A sky130_fd_sc_hd__buf_12
Xfanout1762 _17911_/Q vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__buf_12
Xfanout1773 _12471_/A0 vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__buf_6
XFILLER_38_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19644_ _19644_/CLK _19644_/D vssd1 vssd1 vccd1 vccd1 _19644_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1784 _17905_/Q vssd1 vssd1 vccd1 vccd1 _08874_/D sky130_fd_sc_hd__buf_12
X_16856_ _18745_/Q _12276_/A _16877_/B1 input240/X _12488_/A vssd1 vssd1 vccd1 vccd1
+ _16856_/X sky130_fd_sc_hd__a221o_2
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1795 _17902_/Q vssd1 vssd1 vccd1 vccd1 _12755_/A sky130_fd_sc_hd__buf_4
XFILLER_238_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15807_ _18599_/Q _17697_/A0 _15829_/S vssd1 vssd1 vccd1 vccd1 _18599_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19575_ _19575_/CLK _19575_/D vssd1 vssd1 vccd1 vccd1 _19575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16787_ _16787_/A _16787_/B _16791_/C vssd1 vssd1 vccd1 vccd1 _19283_/D sky130_fd_sc_hd__nor3_1
XFILLER_281_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13999_ _17964_/Q _14032_/B _13998_/Y _14029_/C1 vssd1 vssd1 vccd1 vccd1 _17964_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18526_ _19286_/CLK _18526_/D vssd1 vssd1 vccd1 vccd1 _18526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ _15738_/A _15756_/B vssd1 vssd1 vccd1 vccd1 _15738_/X sky130_fd_sc_hd__xor2_1
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18457_ _19636_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15669_ _19481_/Q _19415_/Q vssd1 vssd1 vccd1 vccd1 _15671_/A sky130_fd_sc_hd__and2_1
XANTENNA_190 _13723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17408_ _18104_/Q _17437_/A2 _17129_/Y _17390_/Y _17407_/X vssd1 vssd1 vccd1 vccd1
+ _17408_/X sky130_fd_sc_hd__a2111o_1
X_09190_ _11452_/A _17702_/A0 _09189_/X vssd1 vssd1 vccd1 vccd1 _11812_/A sky130_fd_sc_hd__o21ai_4
X_18388_ _19465_/CLK _18388_/D vssd1 vssd1 vccd1 vccd1 _18388_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17339_ _19467_/Q _17581_/A _17377_/S vssd1 vssd1 vccd1 vccd1 _17340_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19009_ _19624_/CLK _19009_/D vssd1 vssd1 vccd1 vccd1 _19009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08974_ _11513_/A1 _19110_/Q _19142_/Q _11503_/S0 vssd1 vssd1 vccd1 vccd1 _08974_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_102_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ _18538_/Q _18413_/Q _18022_/Q _17990_/Q _09680_/B1 _10266_/S1 vssd1 vssd1
+ vccd1 vccd1 _09526_/X sky130_fd_sc_hd__mux4_1
XFILLER_213_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _09457_/A _09457_/B vssd1 vssd1 vccd1 vccd1 _09457_/Y sky130_fd_sc_hd__nor2_8
XFILLER_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09388_ _18024_/Q _17992_/Q _10128_/B vssd1 vssd1 vccd1 vccd1 _09388_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ _18640_/Q _18062_/Q _19081_/Q _18985_/Q _11604_/S _11357_/S1 vssd1 vssd1
+ vccd1 vccd1 _11351_/B sky130_fd_sc_hd__mux4_2
XFILLER_193_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10301_ _10297_/X _10300_/X _10301_/S vssd1 vssd1 vccd1 vccd1 _10301_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11281_ _18251_/Q _18826_/Q _18454_/Q _18355_/Q _11284_/B2 _11622_/A1 vssd1 vssd1
+ vccd1 vccd1 _11282_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ input6/X _12552_/X _13013_/X _13019_/X _12538_/B vssd1 vssd1 vccd1 vccd1
+ _13020_/X sky130_fd_sc_hd__o221a_2
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10232_ _11634_/A vssd1 vssd1 vccd1 vccd1 _10232_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1003 _10414_/A2 vssd1 vssd1 vccd1 vccd1 _16486_/A0 sky130_fd_sc_hd__clkbuf_2
X_10163_ _10309_/B _10163_/B vssd1 vssd1 vccd1 vccd1 _10163_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1014 _15047_/Y vssd1 vssd1 vccd1 vccd1 _15076_/S sky130_fd_sc_hd__buf_12
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1025 _16292_/A0 vssd1 vssd1 vccd1 vccd1 _17723_/A0 sky130_fd_sc_hd__buf_6
Xfanout1036 _09491_/X vssd1 vssd1 vccd1 vccd1 _15808_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1047 _17545_/C1 vssd1 vssd1 vccd1 vccd1 _17539_/C1 sky130_fd_sc_hd__buf_4
XFILLER_120_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14971_ _18498_/Q _15011_/A2 _14970_/Y _14991_/C1 vssd1 vssd1 vccd1 vccd1 _18498_/D
+ sky130_fd_sc_hd__a211o_1
X_10094_ _11017_/A1 _19225_/Q _19193_/Q _10168_/S _11397_/A1 vssd1 vssd1 vccd1 vccd1
+ _10094_/X sky130_fd_sc_hd__a221o_1
XFILLER_59_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1058 _15523_/S vssd1 vssd1 vccd1 vccd1 _15498_/S sky130_fd_sc_hd__buf_8
Xfanout1069 _14036_/A vssd1 vssd1 vccd1 vccd1 _14020_/B sky130_fd_sc_hd__clkbuf_4
X_16710_ _19256_/Q _16717_/D _16808_/A vssd1 vssd1 vccd1 vccd1 _16710_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_275_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13922_ _19422_/Q _12579_/Y _12771_/X _13921_/X _12581_/Y vssd1 vssd1 vccd1 vccd1
+ _13922_/X sky130_fd_sc_hd__a221o_1
XFILLER_235_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17690_ _17690_/A0 _19617_/Q _17690_/S vssd1 vssd1 vccd1 vccd1 _19617_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16641_ _16752_/A _16641_/B vssd1 vssd1 vccd1 vccd1 _16641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_207_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13853_ _19388_/Q _13884_/A2 _13851_/X _13852_/X _13884_/C1 vssd1 vssd1 vccd1 vccd1
+ _13853_/X sky130_fd_sc_hd__o221a_4
XFILLER_16_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19360_ _19458_/CLK _19360_/D vssd1 vssd1 vccd1 vccd1 _19360_/Q sky130_fd_sc_hd__dfxtp_1
X_12804_ _12680_/Y _12669_/X _12823_/A vssd1 vssd1 vccd1 vccd1 _12804_/X sky130_fd_sc_hd__mux2_1
X_16572_ _11376_/B _19176_/Q _16586_/S vssd1 vssd1 vccd1 vccd1 _19176_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10996_ _09129_/S _10994_/X _10995_/X _10996_/B1 vssd1 vssd1 vccd1 vccd1 _10996_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_188_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13784_ _19354_/Q _13883_/A2 _13883_/B1 _19482_/Q _13883_/C1 vssd1 vssd1 vccd1 vccd1
+ _13784_/X sky130_fd_sc_hd__a221o_1
XFILLER_215_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18311_ _19634_/CLK _18311_/D vssd1 vssd1 vccd1 vccd1 _18311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ _19474_/Q _15522_/X _15523_/S vssd1 vssd1 vccd1 vccd1 _15523_/X sky130_fd_sc_hd__mux2_1
X_19291_ _19291_/CLK _19291_/D vssd1 vssd1 vccd1 vccd1 _19291_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12821_/A _12821_/B _12734_/Y vssd1 vssd1 vccd1 vccd1 _12735_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18242_ _18817_/CLK _18242_/D vssd1 vssd1 vccd1 vccd1 _18242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _14238_/A _15786_/A2 _15455_/A _15452_/Y vssd1 vssd1 vccd1 vccd1 _15487_/A
+ sky130_fd_sc_hd__o211a_1
X_12666_ _12756_/A _12740_/B vssd1 vssd1 vccd1 vccd1 _12721_/S sky130_fd_sc_hd__nor2_4
XFILLER_169_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14405_ _16314_/A0 _18256_/Q _14416_/S vssd1 vssd1 vccd1 vccd1 _18256_/D sky130_fd_sc_hd__mux2_1
X_11617_ _19098_/Q _19002_/Q _11617_/S vssd1 vssd1 vccd1 vccd1 _11617_/X sky130_fd_sc_hd__mux2_1
X_18173_ _19047_/CLK _18173_/D vssd1 vssd1 vccd1 vccd1 _18173_/Q sky130_fd_sc_hd__dfxtp_1
X_12597_ _12597_/A _12597_/B vssd1 vssd1 vccd1 vccd1 _12597_/Y sky130_fd_sc_hd__nor2_1
X_15385_ _15385_/A _15385_/B vssd1 vssd1 vccd1 vccd1 _15391_/A sky130_fd_sc_hd__and2_1
XFILLER_11_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17124_ _17124_/A _17124_/B _17123_/Y vssd1 vssd1 vccd1 vccd1 _17124_/X sky130_fd_sc_hd__or3b_1
X_14336_ _18193_/Q _17720_/A0 _14338_/S vssd1 vssd1 vccd1 vccd1 _18193_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11548_ _13794_/A _11639_/B _13797_/S vssd1 vssd1 vccd1 vccd1 _11638_/A sky130_fd_sc_hd__a21oi_4
XFILLER_237_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17055_ _19361_/Q _17113_/B vssd1 vssd1 vccd1 vccd1 _17055_/X sky130_fd_sc_hd__or2_1
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14267_ _18305_/Q _14267_/A2 _14266_/X _14442_/B vssd1 vssd1 vccd1 vccd1 _18131_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11479_ _18887_/Q _11479_/B vssd1 vssd1 vccd1 vccd1 _11479_/X sky130_fd_sc_hd__or2_1
X_16006_ _18718_/Q _16016_/A2 _16147_/A2 _18767_/Q _16018_/C1 vssd1 vssd1 vccd1 vccd1
+ _16006_/X sky130_fd_sc_hd__a221o_1
XFILLER_143_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13218_ _13929_/A1 _13217_/X _13204_/X vssd1 vssd1 vccd1 vccd1 _13218_/Y sky130_fd_sc_hd__a21oi_1
X_14198_ _18710_/Q _18097_/Q _14200_/S vssd1 vssd1 vccd1 vccd1 _14199_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13188_/B _13149_/B vssd1 vssd1 vccd1 vccd1 _13149_/X sky130_fd_sc_hd__or2_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17957_ _17958_/CLK _17957_/D vssd1 vssd1 vccd1 vccd1 _17957_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16908_ _16960_/A _16908_/B vssd1 vssd1 vccd1 vccd1 _19311_/D sky130_fd_sc_hd__and2_1
XFILLER_111_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1570 _08897_/Y vssd1 vssd1 vccd1 vccd1 _11508_/B1 sky130_fd_sc_hd__buf_12
Xfanout1581 _08896_/Y vssd1 vssd1 vccd1 vccd1 fanout1581/X sky130_fd_sc_hd__buf_12
X_17888_ _17901_/CLK _17888_/D vssd1 vssd1 vccd1 vccd1 _17888_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1592 _08895_/Y vssd1 vssd1 vccd1 vccd1 _10211_/A1 sky130_fd_sc_hd__buf_12
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19627_ _19627_/CLK _19627_/D vssd1 vssd1 vccd1 vccd1 _19627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16839_ _16839_/A _16839_/B vssd1 vssd1 vccd1 vccd1 _16981_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19558_ _19592_/CLK _19558_/D vssd1 vssd1 vccd1 vccd1 _19558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19159_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09311_ _11503_/S1 _09305_/X _09308_/X _11053_/A vssd1 vssd1 vccd1 vccd1 _09311_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_280_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18509_ _19320_/CLK _18509_/D vssd1 vssd1 vccd1 vccd1 _18509_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19489_ _19525_/CLK _19489_/D vssd1 vssd1 vccd1 vccd1 _19489_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_90_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09242_ input170/X input142/X _09990_/S vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__mux2_4
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09173_ _09166_/X _09172_/X _09163_/X _09169_/X _12466_/A0 _12408_/A vssd1 vssd1
+ vccd1 vccd1 _09173_/X sky130_fd_sc_hd__mux4_2
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput106 dout0[9] vssd1 vssd1 vccd1 vccd1 input106/X sky130_fd_sc_hd__clkbuf_2
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput117 dout1[19] vssd1 vssd1 vccd1 vccd1 input117/X sky130_fd_sc_hd__clkbuf_2
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput128 dout1[29] vssd1 vssd1 vccd1 vccd1 input128/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput139 dout1[39] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_hd__buf_2
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ _08958_/A _08958_/B vssd1 vssd1 vccd1 vccd1 _08957_/Y sky130_fd_sc_hd__nor2_4
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ _11663_/A vssd1 vssd1 vccd1 vccd1 _14346_/B sky130_fd_sc_hd__clkinv_4
XFILLER_263_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _10850_/A1 _17778_/Q _10853_/S _18327_/Q _10557_/S vssd1 vssd1 vccd1 vccd1
+ _10850_/X sky130_fd_sc_hd__o221a_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09509_ _18538_/Q _18413_/Q _09724_/S vssd1 vssd1 vccd1 vccd1 _09509_/X sky130_fd_sc_hd__mux2_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10781_ _11577_/S _10776_/X _10780_/X vssd1 vssd1 vccd1 vccd1 _10781_/Y sky130_fd_sc_hd__o21ai_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12538_/A _12576_/A vssd1 vssd1 vccd1 vccd1 _12580_/A sky130_fd_sc_hd__or2_4
XFILLER_169_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12756_/A _12587_/B vssd1 vssd1 vccd1 vccd1 _12451_/X sky130_fd_sc_hd__and2_1
XFILLER_138_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11402_ _11478_/S _11401_/X _09099_/A vssd1 vssd1 vccd1 vccd1 _11402_/X sky130_fd_sc_hd__a21o_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15170_ _18565_/Q _15351_/A2 _15169_/X _17352_/A vssd1 vssd1 vccd1 vccd1 _18565_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12382_ _12382_/A _12382_/B vssd1 vssd1 vccd1 vccd1 _12382_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_90 _10505_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121_ _17704_/A0 _18060_/Q _14139_/S vssd1 vssd1 vccd1 vccd1 _18060_/D sky130_fd_sc_hd__mux2_1
XFILLER_193_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11333_ _11333_/A1 _11299_/X _11332_/X _11800_/B vssd1 vssd1 vccd1 vccd1 _11828_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ _17669_/A0 _17994_/Q _14072_/S vssd1 vssd1 vccd1 vccd1 _17994_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11264_ _11284_/A1 _18322_/Q _17773_/Q _11284_/B2 vssd1 vssd1 vccd1 vccd1 _11264_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13003_ _13863_/B2 _12998_/X _13002_/X _12704_/S _13000_/Y vssd1 vssd1 vccd1 vccd1
+ _13003_/X sky130_fd_sc_hd__o221a_4
X_10215_ _18623_/Q _18194_/Q _10215_/S vssd1 vssd1 vccd1 vccd1 _10215_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_140_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18860_ _19148_/CLK _18860_/D vssd1 vssd1 vccd1 vccd1 _18860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11195_ _11183_/Y _11187_/Y _11194_/Y vssd1 vssd1 vccd1 vccd1 _11195_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17811_ _19490_/CLK _17811_/D vssd1 vssd1 vccd1 vccd1 _17811_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_267_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10146_ _10143_/X _10144_/X _10145_/X _10297_/A1 _10301_/S vssd1 vssd1 vccd1 vccd1
+ _10146_/X sky130_fd_sc_hd__a221o_1
X_18791_ _19208_/CLK _18791_/D vssd1 vssd1 vccd1 vccd1 _18791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17742_ _18642_/Q vssd1 vssd1 vccd1 vccd1 _18642_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_130_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14954_ _14952_/X _14953_/X _14995_/A1 vssd1 vssd1 vccd1 vccd1 _14954_/X sky130_fd_sc_hd__a21o_1
X_10077_ _09404_/Y _11748_/B _13154_/S vssd1 vssd1 vccd1 vccd1 _11750_/B sky130_fd_sc_hd__o21ai_4
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ _17917_/Q _13971_/A2 _13899_/Y _13903_/X _13579_/A vssd1 vssd1 vccd1 vccd1
+ _13905_/X sky130_fd_sc_hd__a221o_1
XFILLER_236_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17673_ _17706_/A0 _19600_/Q _17690_/S vssd1 vssd1 vccd1 vccd1 _19600_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14885_ _15835_/B _14884_/Y _15006_/B1 vssd1 vssd1 vccd1 vccd1 _14885_/X sky130_fd_sc_hd__a21bo_1
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19412_ _19485_/CLK _19412_/D vssd1 vssd1 vccd1 vccd1 _19412_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_263_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16624_ _19227_/Q input247/X _16627_/S vssd1 vssd1 vccd1 vccd1 _19227_/D sky130_fd_sc_hd__mux2_1
X_13836_ _18128_/Q _13837_/B vssd1 vssd1 vccd1 vccd1 _13900_/C sky130_fd_sc_hd__and2_2
XFILLER_63_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _19471_/CLK _19343_/D vssd1 vssd1 vccd1 vccd1 _19343_/Q sky130_fd_sc_hd__dfxtp_1
X_16555_ _17688_/A0 _19160_/Q _16556_/S vssd1 vssd1 vccd1 vccd1 _19160_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13767_ _12732_/S _13092_/X _13094_/X _13896_/B2 vssd1 vssd1 vccd1 vccd1 _13767_/X
+ sky130_fd_sc_hd__o22a_1
X_10979_ _11365_/B2 _16545_/A0 _10978_/X _11133_/B2 vssd1 vssd1 vccd1 vccd1 _15526_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15506_ _15506_/A _15506_/B vssd1 vssd1 vccd1 vccd1 _15554_/A sky130_fd_sc_hd__xnor2_1
X_19274_ _19276_/CLK _19274_/D vssd1 vssd1 vccd1 vccd1 _19274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12718_ _12710_/X _12717_/X _13041_/S vssd1 vssd1 vccd1 vccd1 _12719_/B sky130_fd_sc_hd__mux2_1
X_16486_ _16486_/A0 _19093_/Q _16488_/S vssd1 vssd1 vccd1 vccd1 _19093_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13698_ _13761_/B _14151_/A vssd1 vssd1 vccd1 vccd1 _13698_/Y sky130_fd_sc_hd__nand2_1
X_18225_ _19226_/CLK _18225_/D vssd1 vssd1 vccd1 vccd1 _18225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15437_ _12788_/B _15436_/X _15437_/B1 vssd1 vssd1 vccd1 vccd1 _15437_/X sky130_fd_sc_hd__a21o_1
X_12649_ _10527_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _12649_/X sky130_fd_sc_hd__and2b_1
XFILLER_50_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18156_ _19644_/CLK _18156_/D vssd1 vssd1 vccd1 vccd1 _18156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15368_ _15456_/A _15368_/B vssd1 vssd1 vccd1 vccd1 _15369_/C sky130_fd_sc_hd__nand2_1
XFILLER_8_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17107_ _19387_/Q _17107_/B vssd1 vssd1 vccd1 vccd1 _17107_/X sky130_fd_sc_hd__or2_1
X_14319_ _18176_/Q _17703_/A0 _14338_/S vssd1 vssd1 vccd1 vccd1 _18176_/D sky130_fd_sc_hd__mux2_1
X_18087_ _18700_/CLK _18087_/D vssd1 vssd1 vccd1 vccd1 _18087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15299_ _15299_/A _15299_/B vssd1 vssd1 vccd1 vccd1 _15299_/Y sky130_fd_sc_hd__xnor2_1
X_17038_ _17202_/B _17046_/A2 _17037_/X _17592_/B vssd1 vssd1 vccd1 vccd1 _19355_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout807 _15817_/S vssd1 vssd1 vccd1 vccd1 _15832_/S sky130_fd_sc_hd__buf_8
XFILLER_98_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09860_ _09859_/A _16462_/A0 _09859_/Y _11800_/B vssd1 vssd1 vccd1 vccd1 _11788_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_113_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout818 _14325_/S vssd1 vssd1 vccd1 vccd1 _14335_/S sky130_fd_sc_hd__buf_12
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout829 _11990_/Y vssd1 vssd1 vccd1 vccd1 _12019_/S sky130_fd_sc_hd__buf_12
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09791_ _10589_/S _09790_/Y _09789_/Y _08874_/D vssd1 vssd1 vccd1 vccd1 _09791_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_274_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18989_ _19636_/CLK _18989_/D vssd1 vssd1 vccd1 vccd1 _18989_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09225_ _11518_/B2 _17702_/A0 _09224_/X _09523_/A vssd1 vssd1 vccd1 vccd1 _15303_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_195_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09156_ _09245_/A _11556_/B _09245_/C _09156_/D vssd1 vssd1 vccd1 vccd1 _09156_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09087_ _11579_/A _12442_/B vssd1 vssd1 vccd1 vccd1 _09087_/Y sky130_fd_sc_hd__nand2_4
XFILLER_190_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ _11157_/A1 _19131_/Q _10001_/S _19099_/Q _11567_/S vssd1 vssd1 vccd1 vccd1
+ _10000_/X sky130_fd_sc_hd__o221a_1
XFILLER_249_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09989_ _09326_/B _09987_/B _09245_/A vssd1 vssd1 vccd1 vccd1 _09989_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ _11953_/B2 _11909_/B _11953_/A2 input239/X vssd1 vssd1 vccd1 vccd1 _11951_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_218_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _10887_/Y _10900_/X _10901_/X vssd1 vssd1 vccd1 vccd1 _10902_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _14671_/A _14680_/C vssd1 vssd1 vccd1 vccd1 _14670_/Y sky130_fd_sc_hd__nor2_2
X_11882_ _11899_/A _11882_/B _11882_/C vssd1 vssd1 vccd1 vccd1 _11882_/X sky130_fd_sc_hd__and3_4
XFILLER_260_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10833_ _09034_/B _09658_/X _09326_/A vssd1 vssd1 vccd1 vccd1 _10834_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13621_ _13614_/Y _13617_/Y _13619_/Y _13620_/X vssd1 vssd1 vccd1 vccd1 _13621_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16340_ _18952_/Q _17672_/A0 _16357_/S vssd1 vssd1 vccd1 vccd1 _18952_/D sky130_fd_sc_hd__mux2_1
XFILLER_260_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13552_ _17874_/Q _13747_/A2 _13550_/X _13682_/B2 vssd1 vssd1 vccd1 vccd1 _13552_/X
+ sky130_fd_sc_hd__a22o_1
X_10764_ _11572_/A1 _19216_/Q _19184_/Q _11325_/S _11584_/C1 vssd1 vssd1 vccd1 vccd1
+ _10764_/X sky130_fd_sc_hd__a221o_1
XFILLER_13_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12503_ _12553_/D _12563_/A vssd1 vssd1 vccd1 vccd1 _12503_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16271_ _16602_/A0 _18885_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _18885_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13483_ _13512_/B _13483_/B vssd1 vssd1 vccd1 vccd1 _13483_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10695_ _18155_/Q _09457_/Y _10694_/X _11406_/B2 vssd1 vssd1 vccd1 vccd1 _10695_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_201_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18010_ _19612_/CLK _18010_/D vssd1 vssd1 vccd1 vccd1 _18010_/Q sky130_fd_sc_hd__dfxtp_1
X_12434_ _15549_/A _12408_/B _12433_/X _13981_/C1 vssd1 vssd1 vccd1 vccd1 _17919_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15222_ _15263_/C _15222_/B vssd1 vssd1 vccd1 vccd1 _15223_/B sky130_fd_sc_hd__xnor2_1
XFILLER_166_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12365_ _17896_/Q _12421_/A _12364_/Y _13981_/C1 vssd1 vssd1 vccd1 vccd1 _17896_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15153_ _18104_/Q _15133_/Y _15152_/X _15216_/A1 vssd1 vssd1 vccd1 vccd1 _15155_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14104_ _16455_/A1 _18044_/Q _14104_/S vssd1 vssd1 vccd1 vccd1 _18044_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11316_ _11314_/X _11315_/X _11577_/S vssd1 vssd1 vccd1 vccd1 _11316_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15084_ _19380_/Q _15092_/B _15084_/C vssd1 vssd1 vccd1 vccd1 _15093_/A sky130_fd_sc_hd__and3_1
XFILLER_126_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12296_ _14688_/B _14675_/A vssd1 vssd1 vccd1 vccd1 _14671_/A sky130_fd_sc_hd__or2_2
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14035_ _12461_/Y _13928_/X _14034_/X _16153_/D vssd1 vssd1 vccd1 vccd1 _17982_/D
+ sky130_fd_sc_hd__o211a_1
X_18912_ _19623_/CLK _18912_/D vssd1 vssd1 vccd1 vccd1 _18912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11247_ _18609_/Q _18180_/Q _11247_/S vssd1 vssd1 vccd1 vccd1 _11247_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18843_ _18875_/CLK _18843_/D vssd1 vssd1 vccd1 vccd1 _18843_/Q sky130_fd_sc_hd__dfxtp_1
X_11178_ _09611_/A _11144_/X _11257_/C1 vssd1 vssd1 vccd1 vccd1 _11178_/X sky130_fd_sc_hd__o21a_1
XFILLER_256_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10129_ _18078_/Q _10364_/B _10128_/X _10346_/S vssd1 vssd1 vccd1 vccd1 _10129_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18774_ _18775_/CLK _18774_/D vssd1 vssd1 vccd1 vccd1 _18774_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ _18708_/Q _16016_/A2 _16004_/B1 _18757_/Q _16004_/C1 vssd1 vssd1 vccd1 vccd1
+ _15986_/X sky130_fd_sc_hd__a221o_1
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17725_ _08991_/A _17724_/B _17724_/Y _17725_/C1 vssd1 vssd1 vccd1 vccd1 _19650_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_264_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14937_ input59/X input94/X _14947_/S vssd1 vssd1 vccd1 vccd1 _14938_/A sky130_fd_sc_hd__mux2_2
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ _17722_/A0 _19584_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _19584_/D sky130_fd_sc_hd__mux2_1
X_14868_ _15009_/A1 _18271_/Q _14867_/Y _14918_/B1 vssd1 vssd1 vccd1 vccd1 _14868_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_24_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16607_ _16607_/A0 _19210_/Q _16618_/S vssd1 vssd1 vccd1 vccd1 _19210_/D sky130_fd_sc_hd__mux2_1
XFILLER_223_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13819_ _17850_/Q _13844_/A2 _13844_/B1 _17882_/Q vssd1 vssd1 vccd1 vccd1 _13819_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17587_ _17587_/A _17589_/B vssd1 vssd1 vccd1 vccd1 _17587_/X sky130_fd_sc_hd__or2_1
XFILLER_250_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14799_ _12459_/X _13996_/B _14683_/X _18637_/Q vssd1 vssd1 vccd1 vccd1 _14799_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_259_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19326_ _19326_/CLK _19326_/D vssd1 vssd1 vccd1 vccd1 _19326_/Q sky130_fd_sc_hd__dfxtp_1
X_16538_ _16538_/A0 _19143_/Q _16556_/S vssd1 vssd1 vccd1 vccd1 _19143_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19257_ _19261_/CLK _19257_/D vssd1 vssd1 vccd1 vccd1 _19257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16469_ _16535_/A0 _19076_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _19076_/D sky130_fd_sc_hd__mux2_1
X_09010_ _18197_/Q _18268_/Q vssd1 vssd1 vccd1 vccd1 _09010_/Y sky130_fd_sc_hd__nand2_2
X_18208_ _19592_/CLK _18208_/D vssd1 vssd1 vccd1 vccd1 _18208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19188_ _19642_/CLK _19188_/D vssd1 vssd1 vccd1 vccd1 _19188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18139_ _19624_/CLK _18139_/D vssd1 vssd1 vccd1 vccd1 _18139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09912_ _18533_/Q _18408_/Q _11481_/C vssd1 vssd1 vccd1 vccd1 _09912_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout604 _17475_/A2 vssd1 vssd1 vccd1 vccd1 _15118_/A sky130_fd_sc_hd__buf_6
Xfanout615 _17558_/B vssd1 vssd1 vccd1 vccd1 _17622_/A2 sky130_fd_sc_hd__buf_4
XFILLER_99_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout626 _16927_/S vssd1 vssd1 vccd1 vccd1 _16967_/S sky130_fd_sc_hd__buf_4
XFILLER_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout637 _17555_/X vssd1 vssd1 vccd1 vccd1 _17589_/B sky130_fd_sc_hd__buf_4
X_09843_ _19069_/Q _18973_/Q _09843_/S vssd1 vssd1 vccd1 vccd1 _09843_/X sky130_fd_sc_hd__mux2_1
Xfanout648 _17077_/B vssd1 vssd1 vccd1 vccd1 _17113_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_98_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout659 _13243_/B1 vssd1 vssd1 vccd1 vccd1 _13781_/B1 sky130_fd_sc_hd__buf_4
XFILLER_274_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09774_ _09768_/Y _09773_/X _11332_/B1 vssd1 vssd1 vccd1 vccd1 _11790_/D sky130_fd_sc_hd__a21oi_4
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09208_ _09196_/X _09207_/X _10301_/S vssd1 vssd1 vccd1 vccd1 _09208_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10480_ _11566_/A1 _18229_/Q _10840_/S _18964_/Q vssd1 vssd1 vccd1 vccd1 _10480_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_183_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09139_ _11024_/A1 _09138_/X _11257_/C1 _09105_/X vssd1 vssd1 vccd1 vccd1 _09139_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_185_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12150_ _17845_/Q _12152_/C _12149_/Y vssd1 vssd1 vccd1 vccd1 _17845_/D sky130_fd_sc_hd__o21a_1
XFILLER_151_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11101_ _10532_/A _11067_/X _11800_/B vssd1 vssd1 vccd1 vccd1 _11101_/X sky130_fd_sc_hd__o21a_1
XFILLER_190_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12081_ _17818_/Q _12087_/B vssd1 vssd1 vccd1 vccd1 _12081_/X sky130_fd_sc_hd__or2_1
XFILLER_2_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11032_ _11428_/A _11031_/X _11501_/B1 vssd1 vssd1 vccd1 vccd1 _11032_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _15843_/A _15840_/B vssd1 vssd1 vccd1 vccd1 _15840_/Y sky130_fd_sc_hd__nand2_1
XFILLER_265_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _18592_/Q _15772_/B vssd1 vssd1 vccd1 vccd1 _15791_/B sky130_fd_sc_hd__nand2_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12983_ _13421_/A _11737_/X _12982_/Y _09866_/B vssd1 vssd1 vccd1 vccd1 _12983_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _11643_/Y _17520_/A2 _17532_/A2 _17814_/Q _17538_/A vssd1 vssd1 vccd1 vccd1
+ _17510_/X sky130_fd_sc_hd__a221o_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _18629_/Q _14683_/A _14683_/B _14912_/A1 _12922_/Y vssd1 vssd1 vccd1 vccd1
+ _14722_/X sky130_fd_sc_hd__a32o_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18490_ _19286_/CLK _18490_/D vssd1 vssd1 vccd1 vccd1 _18490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _11939_/A1 _11831_/B _11949_/B1 input220/X vssd1 vssd1 vccd1 vccd1 _11934_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_520 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_531 _18573_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_542 _18104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_178_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18741_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17441_ _18572_/Q _15103_/Y _17546_/A2 vssd1 vssd1 vccd1 vccd1 _17441_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14653_ _16314_/A0 _18459_/Q _14664_/S vssd1 vssd1 vccd1 vccd1 _18459_/D sky130_fd_sc_hd__mux2_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _11865_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11865_/Y sky130_fd_sc_hd__nand2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19306_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13604_ _13791_/A _13595_/Y _13596_/X _13611_/B _13622_/A vssd1 vssd1 vccd1 vccd1
+ _13604_/X sky130_fd_sc_hd__a32o_1
XFILLER_220_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10816_ _18896_/Q _10816_/A2 _08899_/A vssd1 vssd1 vccd1 vccd1 _10816_/X sky130_fd_sc_hd__o21a_1
X_17372_ _17592_/B _17372_/B vssd1 vssd1 vccd1 vccd1 _19483_/D sky130_fd_sc_hd__and2_1
X_11796_ _11816_/A _11796_/B vssd1 vssd1 vccd1 vccd1 _11825_/B sky130_fd_sc_hd__nor2_8
X_14584_ _14592_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _18400_/D sky130_fd_sc_hd__or2_1
X_19111_ _19157_/CLK _19111_/D vssd1 vssd1 vccd1 vccd1 _19111_/Q sky130_fd_sc_hd__dfxtp_1
X_16323_ _17721_/A0 _18936_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _18936_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ _13797_/A0 _12756_/Y _13535_/S vssd1 vssd1 vccd1 vccd1 _13535_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ _10747_/A1 _10746_/X _08898_/Y vssd1 vssd1 vccd1 vccd1 _10747_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19042_ _19625_/CLK _19042_/D vssd1 vssd1 vccd1 vccd1 _19042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16254_ _17718_/A0 _18869_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _18869_/D sky130_fd_sc_hd__mux2_1
X_10678_ _09034_/B _09487_/X _09326_/A vssd1 vssd1 vccd1 vccd1 _10679_/B sky130_fd_sc_hd__a21oi_2
XFILLER_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13466_ _13466_/A _13466_/B vssd1 vssd1 vccd1 vccd1 _14145_/B sky130_fd_sc_hd__nor2_1
XFILLER_174_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15205_ _19461_/Q _15204_/Y _15400_/S vssd1 vssd1 vccd1 vccd1 _15205_/X sky130_fd_sc_hd__mux2_1
X_12417_ _12429_/A1 _09232_/A _09146_/X _12417_/B1 _18399_/Q vssd1 vssd1 vccd1 vccd1
+ _12418_/B sky130_fd_sc_hd__o32ai_2
X_16185_ _16615_/A0 _18802_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _18802_/D sky130_fd_sc_hd__mux2_1
XFILLER_182_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13397_ _18115_/Q _18114_/Q _13397_/C vssd1 vssd1 vccd1 vccd1 _13406_/B sky130_fd_sc_hd__and3_1
XFILLER_160_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15136_ _15137_/A _15137_/B vssd1 vssd1 vccd1 vccd1 _15138_/B sky130_fd_sc_hd__nor2_1
X_12348_ _12420_/A1 _09907_/A _09738_/X _12420_/B1 _18376_/Q vssd1 vssd1 vccd1 vccd1
+ _12349_/B sky130_fd_sc_hd__o32ai_4
XFILLER_142_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12279_ _18093_/Q _12305_/A2 _12305_/B1 _18516_/Q vssd1 vssd1 vccd1 vccd1 _12483_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_141_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15067_ _18551_/Q _17711_/A0 _15079_/S vssd1 vssd1 vccd1 vccd1 _18551_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ _17974_/Q _14020_/B vssd1 vssd1 vccd1 vccd1 _14018_/X sky130_fd_sc_hd__or2_1
XFILLER_141_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18826_ _19589_/CLK _18826_/D vssd1 vssd1 vccd1 vccd1 _18826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18757_ _18775_/CLK _18757_/D vssd1 vssd1 vccd1 vccd1 _18757_/Q sky130_fd_sc_hd__dfxtp_1
X_15969_ _18700_/Q _15977_/A2 _15968_/X _14177_/A vssd1 vssd1 vccd1 vccd1 _18700_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17708_ _17708_/A0 _19634_/Q _17719_/S vssd1 vssd1 vccd1 vccd1 _19634_/D sky130_fd_sc_hd__mux2_1
X_09490_ _11556_/C _09478_/X _09489_/X _11687_/A vssd1 vssd1 vccd1 vccd1 _09490_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18688_ _19276_/CLK _18688_/D vssd1 vssd1 vccd1 vccd1 _18688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17639_ _17672_/A0 _19567_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _19567_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19309_ _19310_/CLK _19309_/D vssd1 vssd1 vccd1 vccd1 _19309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09826_ _18342_/Q _11224_/B vssd1 vssd1 vccd1 vccd1 _09826_/X sky130_fd_sc_hd__or2_1
XFILLER_101_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout489 _15010_/B1 vssd1 vssd1 vccd1 vccd1 _14950_/B1 sky130_fd_sc_hd__buf_12
XFILLER_219_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09757_ _11565_/A1 _17761_/Q _11073_/B1 _18310_/Q vssd1 vssd1 vccd1 vccd1 _09757_/X
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_5_wb_clk_i _19652_/A vssd1 vssd1 vccd1 vccd1 _19226_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _19622_/Q _18911_/Q _09688_/S vssd1 vssd1 vccd1 vccd1 _09688_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_200_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19055_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_214_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11651_/B _11650_/B vssd1 vssd1 vccd1 vccd1 _11846_/A sky130_fd_sc_hd__or2_4
XFILLER_242_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10601_ _10602_/A _12650_/B vssd1 vssd1 vccd1 vccd1 _10603_/A sky130_fd_sc_hd__and2_4
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11581_ _19066_/Q _19034_/Q _11581_/S vssd1 vssd1 vccd1 vccd1 _11581_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10532_ _10532_/A _10532_/B vssd1 vssd1 vccd1 vccd1 _10532_/Y sky130_fd_sc_hd__nor2_1
X_13320_ _13259_/X _13310_/X _13312_/Y _13319_/X vssd1 vssd1 vccd1 vccd1 _13320_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_210_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13251_ _13928_/A1 _13239_/X _13250_/X vssd1 vssd1 vccd1 vccd1 _13251_/X sky130_fd_sc_hd__a21o_4
X_10463_ _19060_/Q _19028_/Q _10467_/S vssd1 vssd1 vccd1 vccd1 _10463_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12202_ _17865_/Q _12202_/B vssd1 vssd1 vccd1 vccd1 _12208_/C sky130_fd_sc_hd__and2_2
XFILLER_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13182_ _13757_/A _13990_/B _13163_/Y vssd1 vssd1 vccd1 vccd1 _13182_/Y sky130_fd_sc_hd__o21ai_1
X_10394_ _10392_/X _10393_/X _11577_/S vssd1 vssd1 vccd1 vccd1 _10394_/X sky130_fd_sc_hd__mux2_1
X_12133_ _17839_/Q _12136_/C _12219_/A vssd1 vssd1 vccd1 vccd1 _12133_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_151_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17990_ _18445_/CLK _17990_/D vssd1 vssd1 vccd1 vccd1 _17990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1900 _16740_/A vssd1 vssd1 vccd1 vccd1 _16776_/A sky130_fd_sc_hd__buf_2
X_16941_ _18766_/Q _16965_/A2 _16965_/B1 input231/X _16965_/C1 vssd1 vssd1 vccd1 vccd1
+ _16941_/X sky130_fd_sc_hd__a221o_2
X_12064_ _12962_/A0 _12086_/A2 _12063_/X _14342_/A vssd1 vssd1 vccd1 vccd1 _17809_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11015_ _11478_/S _11014_/X _10243_/A vssd1 vssd1 vccd1 vccd1 _11015_/X sky130_fd_sc_hd__a21o_1
XFILLER_238_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16872_ _16928_/A _16872_/B vssd1 vssd1 vccd1 vccd1 _19302_/D sky130_fd_sc_hd__and2_1
XFILLER_277_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18611_ _18613_/CLK _18611_/D vssd1 vssd1 vccd1 vccd1 _18611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout990 _11647_/X vssd1 vssd1 vccd1 vccd1 _11864_/B sky130_fd_sc_hd__clkbuf_8
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ _18615_/Q _17713_/A0 _15833_/S vssd1 vssd1 vccd1 vccd1 _18615_/D sky130_fd_sc_hd__mux2_1
X_19591_ _19591_/CLK _19591_/D vssd1 vssd1 vccd1 vccd1 _19591_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18542_ _19564_/CLK _18542_/D vssd1 vssd1 vccd1 vccd1 _18542_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _19485_/Q _19419_/Q vssd1 vssd1 vccd1 vccd1 _15755_/B sky130_fd_sc_hd__nand2_1
X_12966_ _17827_/Q _13944_/B vssd1 vssd1 vccd1 vccd1 _12966_/X sky130_fd_sc_hd__or2_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _14964_/B1 _14703_/X _14704_/X _14690_/Y vssd1 vssd1 vccd1 vccd1 _14705_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_205_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18473_ _19229_/CLK _18473_/D vssd1 vssd1 vccd1 vccd1 _18473_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11917_ _18571_/Q _11918_/A2 _11706_/B _11751_/Y vssd1 vssd1 vccd1 vccd1 _11917_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_233_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15685_ _15685_/A vssd1 vssd1 vccd1 vccd1 _15689_/A sky130_fd_sc_hd__inv_2
XFILLER_73_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 _10301_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12897_ _13194_/S _12896_/Y _13197_/B1 vssd1 vssd1 vccd1 vccd1 _12897_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_361 _15129_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_372 _18274_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17424_ _19496_/Q _17453_/B _17422_/X _17423_/Y _17328_/A vssd1 vssd1 vccd1 vccd1
+ _19496_/D sky130_fd_sc_hd__o221a_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_383 _15955_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14636_ _17695_/A0 _18442_/Q _14648_/S vssd1 vssd1 vccd1 vccd1 _18442_/D sky130_fd_sc_hd__mux2_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11848_ _11952_/A2 _11845_/X _11847_/X vssd1 vssd1 vccd1 vccd1 _11849_/B sky130_fd_sc_hd__a21oi_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_394 _15082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _19475_/Q _17178_/B _17379_/S vssd1 vssd1 vccd1 vccd1 _17356_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14567_ _18392_/Q _14575_/A2 _14575_/B1 input20/X vssd1 vssd1 vccd1 vccd1 _14568_/B
+ sky130_fd_sc_hd__o22a_1
X_11779_ _11810_/A _11779_/B vssd1 vssd1 vccd1 vccd1 _11779_/X sky130_fd_sc_hd__or2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16306_ _17704_/A0 _18919_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _18919_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13518_ _19250_/Q _13625_/A2 _13625_/B1 _19282_/Q vssd1 vssd1 vccd1 vccd1 _13518_/X
+ sky130_fd_sc_hd__a22o_2
X_17286_ _19446_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17286_/Y sky130_fd_sc_hd__nand2_1
X_14498_ _17700_/A0 _18348_/Q _14517_/S vssd1 vssd1 vccd1 vccd1 _18348_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19025_ _19025_/CLK _19025_/D vssd1 vssd1 vccd1 vccd1 _19025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ _17668_/A0 _18852_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _18852_/D sky130_fd_sc_hd__mux2_1
X_13449_ _17839_/Q _13846_/B vssd1 vssd1 vccd1 vccd1 _13449_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_75_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19595_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_173_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16168_ _17698_/A0 _18785_/Q _16189_/S vssd1 vssd1 vccd1 vccd1 _18785_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15119_ _08882_/B _17445_/C1 _17556_/A vssd1 vssd1 vccd1 vccd1 _15119_/Y sky130_fd_sc_hd__o21ai_2
X_16099_ _18752_/Q _16141_/B vssd1 vssd1 vccd1 vccd1 _16099_/Y sky130_fd_sc_hd__nand2_1
X_08990_ _12053_/A _12051_/A _08932_/A vssd1 vssd1 vccd1 vccd1 _08990_/X sky130_fd_sc_hd__o21ba_2
XFILLER_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09611_ _09611_/A _09611_/B vssd1 vssd1 vccd1 vccd1 _09611_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18809_ _19628_/CLK _18809_/D vssd1 vssd1 vccd1 vccd1 _18809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09542_ _18600_/Q _18171_/Q _09542_/S vssd1 vssd1 vccd1 vccd1 _09542_/X sky130_fd_sc_hd__mux2_1
XFILLER_225_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09473_ _17915_/Q _09643_/A _09472_/X _09367_/B vssd1 vssd1 vccd1 vccd1 _09475_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_252_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1207 _12667_/X vssd1 vssd1 vccd1 vccd1 _12732_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_160_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1218 _12441_/Y vssd1 vssd1 vccd1 vccd1 _12442_/D sky130_fd_sc_hd__buf_4
Xfanout1229 _15329_/B vssd1 vssd1 vccd1 vccd1 _12318_/A sky130_fd_sc_hd__buf_6
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09809_ _11282_/A _09801_/X _09800_/X _11285_/S vssd1 vssd1 vccd1 vccd1 _09809_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_207_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12820_ _12818_/X _12933_/B _12933_/A vssd1 vssd1 vccd1 vccd1 _12820_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _13414_/A _12750_/X _12745_/X vssd1 vssd1 vccd1 vccd1 _12751_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_199_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _14347_/B _11668_/Y _11686_/X _14268_/B _11701_/X vssd1 vssd1 vccd1 vccd1
+ _11702_/X sky130_fd_sc_hd__o32a_4
XFILLER_231_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _19472_/Q _19406_/Q vssd1 vssd1 vccd1 vccd1 _15472_/A sky130_fd_sc_hd__nand2_1
X_12682_ _12681_/X _12680_/A _12821_/A vssd1 vssd1 vccd1 vccd1 _12872_/B sky130_fd_sc_hd__mux2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14421_ _19230_/Q _15014_/B _18274_/D vssd1 vssd1 vccd1 vccd1 _18272_/D sky130_fd_sc_hd__and3_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11634_/A _11634_/B vssd1 vssd1 vccd1 vccd1 _11633_/Y sky130_fd_sc_hd__nor2_1
XFILLER_230_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _19398_/Q fanout534/X _17423_/A _17158_/B2 vssd1 vssd1 vccd1 vccd1 _17141_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_129_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14352_ _18204_/Q _16526_/A0 _14383_/S vssd1 vssd1 vccd1 vccd1 _18204_/D sky130_fd_sc_hd__mux2_1
X_11564_ _11084_/S _11559_/X _11563_/X vssd1 vssd1 vccd1 vccd1 _11564_/X sky130_fd_sc_hd__o21a_1
XFILLER_155_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13303_ input267/X _12575_/Y _13297_/X _13303_/B2 vssd1 vssd1 vccd1 vccd1 _13303_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10515_ _18464_/Q _18365_/Q _10582_/S vssd1 vssd1 vccd1 vccd1 _10515_/X sky130_fd_sc_hd__mux2_1
X_17071_ _19369_/Q _17107_/B vssd1 vssd1 vccd1 vccd1 _17071_/X sky130_fd_sc_hd__or2_1
X_11495_ _11428_/A _11494_/X _11495_/B1 vssd1 vssd1 vccd1 vccd1 _11495_/X sky130_fd_sc_hd__a21o_1
X_14283_ _17701_/A0 _18142_/Q _14304_/S vssd1 vssd1 vccd1 vccd1 _18142_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16022_ _18733_/Q _15854_/A _16034_/S vssd1 vssd1 vccd1 vccd1 _16022_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10446_ _11601_/A _10445_/Y _10444_/Y _11602_/C1 vssd1 vssd1 vccd1 vccd1 _10446_/X
+ sky130_fd_sc_hd__a211o_1
X_13234_ _13227_/X _13231_/Y _13233_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _13234_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ _19304_/Q _13165_/B _13165_/C vssd1 vssd1 vccd1 vccd1 _13165_/X sky130_fd_sc_hd__or3_2
XFILLER_151_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10377_ _13818_/A vssd1 vssd1 vccd1 vccd1 _10377_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12116_ _17832_/Q _12114_/B _12115_/Y vssd1 vssd1 vccd1 vccd1 _17832_/D sky130_fd_sc_hd__o21a_1
XFILLER_3_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17973_ _17975_/CLK _17973_/D vssd1 vssd1 vccd1 vccd1 _17973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13096_ _13896_/B2 _13092_/X _13094_/X _12732_/S _13095_/Y vssd1 vssd1 vccd1 vccd1
+ _13096_/X sky130_fd_sc_hd__o221a_4
XFILLER_285_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1730 _18660_/Q vssd1 vssd1 vccd1 vccd1 _08828_/A sky130_fd_sc_hd__buf_6
X_16924_ _16928_/A _16924_/B vssd1 vssd1 vccd1 vccd1 _19315_/D sky130_fd_sc_hd__and2_1
X_12047_ _17801_/Q _12051_/B vssd1 vssd1 vccd1 vccd1 _12047_/X sky130_fd_sc_hd__or2_1
XFILLER_266_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1741 _18273_/Q vssd1 vssd1 vccd1 vccd1 _14784_/S sky130_fd_sc_hd__buf_12
XFILLER_242_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1752 _17918_/Q vssd1 vssd1 vccd1 vccd1 _12442_/A sky130_fd_sc_hd__buf_12
XFILLER_93_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1763 _12320_/A vssd1 vssd1 vccd1 vccd1 _11579_/A sky130_fd_sc_hd__buf_12
Xfanout1774 _12471_/A0 vssd1 vssd1 vccd1 vccd1 _11481_/A sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_193_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19641_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_266_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1785 _08896_/A vssd1 vssd1 vccd1 vccd1 _10747_/A1 sky130_fd_sc_hd__buf_12
X_16855_ _16928_/A _16855_/B vssd1 vssd1 vccd1 vccd1 _19298_/D sky130_fd_sc_hd__and2_1
X_19643_ _19643_/CLK _19643_/D vssd1 vssd1 vccd1 vccd1 _19643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1796 _08816_/A vssd1 vssd1 vccd1 vccd1 _08932_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_281_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_122_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19324_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15806_ _18598_/Q _16431_/A1 _15829_/S vssd1 vssd1 vccd1 vccd1 _18598_/D sky130_fd_sc_hd__mux2_1
X_19574_ _19649_/CLK _19574_/D vssd1 vssd1 vccd1 vccd1 _19574_/Q sky130_fd_sc_hd__dfxtp_1
X_16786_ _19283_/Q _16786_/B vssd1 vssd1 vccd1 vccd1 _16791_/C sky130_fd_sc_hd__and2_2
X_13998_ _14032_/B _13998_/B vssd1 vssd1 vccd1 vccd1 _13998_/Y sky130_fd_sc_hd__nand2_1
XFILLER_207_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18525_ _19286_/CLK _18525_/D vssd1 vssd1 vccd1 vccd1 _18525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15737_ _15713_/A _15715_/B _15713_/B vssd1 vssd1 vccd1 vccd1 _15756_/B sky130_fd_sc_hd__a21boi_2
XFILLER_240_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12949_ _11734_/B _13230_/A1 _12948_/X _11734_/A vssd1 vssd1 vccd1 vccd1 _12949_/X
+ sky130_fd_sc_hd__o2bb2a_2
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18456_ _19637_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_1
X_15668_ _15651_/B _15653_/B _15651_/A vssd1 vssd1 vccd1 vccd1 _15672_/A sky130_fd_sc_hd__a21bo_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_180 _13527_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_191 _13741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17407_ _18565_/Q _17461_/A2 _17406_/X _17426_/B1 vssd1 vssd1 vccd1 vccd1 _17407_/X
+ sky130_fd_sc_hd__o211a_1
X_14619_ _17711_/A0 _18426_/Q _14631_/S vssd1 vssd1 vccd1 vccd1 _18426_/D sky130_fd_sc_hd__mux2_1
X_18387_ _19466_/CLK _18387_/D vssd1 vssd1 vccd1 vccd1 _18387_/Q sky130_fd_sc_hd__dfxtp_4
X_15599_ _15638_/C vssd1 vssd1 vccd1 vccd1 _15599_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17338_ _17338_/A _17338_/B vssd1 vssd1 vccd1 vccd1 _19466_/D sky130_fd_sc_hd__and2_1
XFILLER_147_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17269_ _14238_/A _17540_/B1 _17473_/A _17313_/B vssd1 vssd1 vccd1 vccd1 _17269_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_19008_ _19653_/A _19008_/D vssd1 vssd1 vccd1 vccd1 _19008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08973_ _11513_/A1 _18950_/Q _18215_/Q _11503_/S0 vssd1 vssd1 vccd1 vccd1 _08973_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ _09948_/B _15214_/A _09476_/X vssd1 vssd1 vccd1 vccd1 _12613_/B sky130_fd_sc_hd__a21boi_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09456_ _10253_/A _19170_/Q _09464_/S vssd1 vssd1 vccd1 vccd1 _09456_/X sky130_fd_sc_hd__and3_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09387_ _10219_/A1 _19562_/Q _10128_/B _19594_/Q _10225_/S vssd1 vssd1 vccd1 vccd1
+ _09387_/X sky130_fd_sc_hd__o221a_1
XFILLER_212_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10300_ _10298_/X _10299_/X _10300_/S vssd1 vssd1 vccd1 vccd1 _10300_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11280_ _11280_/A _11280_/B vssd1 vssd1 vccd1 vccd1 _11280_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10231_ _10233_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__nor2_2
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10162_ _11218_/A _10162_/B vssd1 vssd1 vccd1 vccd1 _10163_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1004 _10385_/X vssd1 vssd1 vccd1 vccd1 _10414_/A2 sky130_fd_sc_hd__buf_12
Xoutput390 _11942_/X vssd1 vssd1 vccd1 vccd1 din0[22] sky130_fd_sc_hd__buf_4
Xfanout1015 _14402_/S vssd1 vssd1 vccd1 vccd1 _14416_/S sky130_fd_sc_hd__buf_12
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1026 _11558_/X vssd1 vssd1 vccd1 vccd1 _16292_/A0 sky130_fd_sc_hd__buf_8
X_10093_ _10243_/A _10093_/B vssd1 vssd1 vccd1 vccd1 _10093_/Y sky130_fd_sc_hd__nor2_1
Xfanout1037 _17698_/A0 vssd1 vssd1 vccd1 vccd1 _17665_/A0 sky130_fd_sc_hd__clkbuf_4
X_14970_ _14966_/Y _14969_/X _15010_/B1 vssd1 vssd1 vccd1 vccd1 _14970_/Y sky130_fd_sc_hd__a21oi_4
Xfanout1048 _17528_/B vssd1 vssd1 vccd1 vccd1 _17545_/C1 sky130_fd_sc_hd__buf_4
XFILLER_102_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1059 _13322_/Y vssd1 vssd1 vccd1 vccd1 _13968_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13921_ _19552_/Q _19520_/Q _13921_/S vssd1 vssd1 vccd1 vccd1 _13921_/X sky130_fd_sc_hd__mux2_1
XFILLER_235_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16640_ _19236_/Q _16643_/C vssd1 vssd1 vccd1 vccd1 _16641_/B sky130_fd_sc_hd__and2_1
XFILLER_75_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13852_ _19356_/Q _13883_/A2 _13883_/B1 _19484_/Q _13883_/C1 vssd1 vssd1 vccd1 vccd1
+ _13852_/X sky130_fd_sc_hd__a221o_1
XFILLER_63_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ _12803_/A vssd1 vssd1 vccd1 vccd1 _12803_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16571_ _11452_/B _19175_/Q _16586_/S vssd1 vssd1 vccd1 vccd1 _19175_/D sky130_fd_sc_hd__mux2_1
X_13783_ _19450_/Q _13949_/A2 _13781_/X _13782_/X _13949_/C1 vssd1 vssd1 vccd1 vccd1
+ _13783_/X sky130_fd_sc_hd__o221a_1
X_10995_ _11469_/A1 _19149_/Q _11386_/S _19117_/Q _10403_/S vssd1 vssd1 vccd1 vccd1
+ _10995_/X sky130_fd_sc_hd__o221a_1
XFILLER_16_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18310_ _19148_/CLK _18310_/D vssd1 vssd1 vccd1 vccd1 _18310_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ _15522_/A _15522_/B vssd1 vssd1 vccd1 vccd1 _15522_/X sky130_fd_sc_hd__xor2_1
X_19290_ _19291_/CLK _19290_/D vssd1 vssd1 vccd1 vccd1 _19290_/Q sky130_fd_sc_hd__dfxtp_1
X_12734_ _12823_/A _12734_/B vssd1 vssd1 vccd1 vccd1 _12734_/Y sky130_fd_sc_hd__nor2_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18241_ _18880_/CLK _18241_/D vssd1 vssd1 vccd1 vccd1 _18241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _14238_/A _15786_/A2 _15452_/Y vssd1 vssd1 vccd1 vccd1 _15455_/B sky130_fd_sc_hd__o21a_1
XFILLER_176_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12665_ _12665_/A _12665_/B _14156_/S vssd1 vssd1 vccd1 vccd1 _12665_/X sky130_fd_sc_hd__or3_1
XFILLER_231_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14404_ _17678_/A0 _18255_/Q _14416_/S vssd1 vssd1 vccd1 vccd1 _18255_/D sky130_fd_sc_hd__mux2_1
X_18172_ _18880_/CLK _18172_/D vssd1 vssd1 vccd1 vccd1 _18172_/Q sky130_fd_sc_hd__dfxtp_1
X_11616_ _11614_/X _11615_/X _11616_/S vssd1 vssd1 vccd1 vccd1 _11616_/X sky130_fd_sc_hd__mux2_1
X_15384_ _15387_/A _15387_/B vssd1 vssd1 vccd1 vccd1 _15384_/Y sky130_fd_sc_hd__nor2_1
X_12596_ _12596_/A _12596_/B vssd1 vssd1 vccd1 vccd1 _12596_/Y sky130_fd_sc_hd__nor2_2
XFILLER_156_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17123_ _17157_/A _17123_/B vssd1 vssd1 vccd1 vccd1 _17123_/Y sky130_fd_sc_hd__nand2_1
X_14335_ _18192_/Q _17719_/A0 _14335_/S vssd1 vssd1 vccd1 vccd1 _18192_/D sky130_fd_sc_hd__mux2_1
X_11547_ _13727_/A _11642_/B _12647_/B _11544_/X vssd1 vssd1 vccd1 vccd1 _11639_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17054_ _17117_/B _17114_/A2 _17053_/X _17378_/A vssd1 vssd1 vccd1 vccd1 _19360_/D
+ sky130_fd_sc_hd__o211a_1
X_14266_ _18131_/Q _14266_/B vssd1 vssd1 vccd1 vccd1 _14266_/X sky130_fd_sc_hd__or2_1
X_11478_ _11476_/X _11477_/X _11478_/S vssd1 vssd1 vccd1 vccd1 _11478_/X sky130_fd_sc_hd__mux2_2
XFILLER_171_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16005_ _18718_/Q _16005_/A2 _16004_/X _14197_/A vssd1 vssd1 vccd1 vccd1 _18718_/D
+ sky130_fd_sc_hd__o211a_1
X_13217_ _13945_/B2 _13205_/X _13216_/X vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__a21o_4
X_10429_ _10419_/S _10421_/X _10420_/X _11507_/S vssd1 vssd1 vccd1 vccd1 _10429_/X
+ sky130_fd_sc_hd__a211o_1
X_14197_ _14197_/A _14197_/B vssd1 vssd1 vccd1 vccd1 _18096_/D sky130_fd_sc_hd__and2_1
XFILLER_98_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _13148_/A _13148_/B _13148_/C vssd1 vssd1 vccd1 vccd1 _13149_/B sky130_fd_sc_hd__and3_1
XFILLER_285_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17956_ _17975_/CLK _17956_/D vssd1 vssd1 vccd1 vccd1 _17956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13079_ _13079_/A _13079_/B _13079_/C vssd1 vssd1 vccd1 vccd1 _13079_/X sky130_fd_sc_hd__and3_1
XFILLER_257_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1560 _08899_/Y vssd1 vssd1 vccd1 vccd1 _09381_/S sky130_fd_sc_hd__buf_8
XFILLER_66_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16907_ _19311_/Q _17589_/A _16963_/S vssd1 vssd1 vccd1 vccd1 _16908_/B sky130_fd_sc_hd__mux2_1
XFILLER_238_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17887_ _19650_/CLK _17887_/D vssd1 vssd1 vccd1 vccd1 _17887_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1571 _11127_/S vssd1 vssd1 vccd1 vccd1 _11361_/S sky130_fd_sc_hd__buf_8
XFILLER_239_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1582 _10881_/S1 vssd1 vssd1 vccd1 vccd1 _11357_/S1 sky130_fd_sc_hd__buf_8
Xfanout1593 _08894_/Y vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__buf_12
XFILLER_65_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19626_ _19626_/CLK _19626_/D vssd1 vssd1 vccd1 vccd1 _19626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_265_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16838_ _17051_/A _16975_/B _17051_/D _17052_/C vssd1 vssd1 vccd1 vccd1 _16843_/C
+ sky130_fd_sc_hd__and4bb_1
XFILLER_281_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16769_ _19277_/Q _16770_/B vssd1 vssd1 vccd1 vccd1 _16771_/B sky130_fd_sc_hd__nor2_1
X_19557_ _19589_/CLK _19557_/D vssd1 vssd1 vccd1 vccd1 _19557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09310_ _11503_/S1 _09300_/X _09309_/X _11438_/B1 vssd1 vssd1 vccd1 vccd1 _09310_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_206_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18508_ _19229_/CLK _18508_/D vssd1 vssd1 vccd1 vccd1 _18508_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19488_ _19525_/CLK _19488_/D vssd1 vssd1 vccd1 vccd1 _19488_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09241_ _09019_/Y _09239_/X _09240_/X vssd1 vssd1 vccd1 vccd1 _09241_/Y sky130_fd_sc_hd__a21oi_1
X_18439_ _19618_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_90_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18749_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09172_ _10169_/S _09170_/X _09171_/X vssd1 vssd1 vccd1 vccd1 _09172_/X sky130_fd_sc_hd__a21o_1
XFILLER_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput107 dout1[0] vssd1 vssd1 vccd1 vccd1 input107/X sky130_fd_sc_hd__clkbuf_2
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput118 dout1[1] vssd1 vssd1 vccd1 vccd1 input118/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08956_ _09055_/B _08956_/B _08956_/C _08956_/D vssd1 vssd1 vccd1 vccd1 _08958_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput129 dout1[2] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08887_ _18590_/Q _11724_/B _08887_/C vssd1 vssd1 vccd1 vccd1 _08887_/Y sky130_fd_sc_hd__nor3_4
XFILLER_111_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09508_ _18313_/Q _17764_/Q _09724_/S vssd1 vssd1 vccd1 vccd1 _09508_/X sky130_fd_sc_hd__mux2_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10785_/A _10779_/X _11563_/B1 vssd1 vssd1 vccd1 vccd1 _10780_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09439_ _19074_/Q _09671_/S _09438_/X _10266_/S1 vssd1 vssd1 vccd1 vccd1 _09439_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12450_ _13421_/A _13462_/A _15083_/A _12461_/A vssd1 vssd1 vccd1 vccd1 _12450_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ _11469_/A1 _18607_/Q _18178_/Q _11477_/S vssd1 vssd1 vccd1 vccd1 _11401_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12381_ _18387_/Q _12429_/B1 _09481_/B _08858_/A vssd1 vssd1 vccd1 vccd1 _12382_/B
+ sky130_fd_sc_hd__a2bb2o_2
XANTENNA_80 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_91 _11864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ _16471_/A0 _18059_/Q _14139_/S vssd1 vssd1 vccd1 vccd1 _18059_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11332_ _11330_/X _11331_/X _11332_/B1 vssd1 vssd1 vccd1 vccd1 _11332_/X sky130_fd_sc_hd__a21o_4
XFILLER_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14051_ _16535_/A0 _17993_/Q _14072_/S vssd1 vssd1 vccd1 vccd1 _17993_/D sky130_fd_sc_hd__mux2_1
XFILLER_193_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11263_ _11277_/A1 _19601_/Q _19569_/Q _11284_/B2 vssd1 vssd1 vccd1 vccd1 _11263_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13002_ _13315_/S _13001_/Y _13413_/B1 vssd1 vssd1 vccd1 vccd1 _13002_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10214_ _18265_/Q _18840_/Q _10215_/S vssd1 vssd1 vccd1 vccd1 _10214_/X sky130_fd_sc_hd__mux2_1
X_11194_ _11194_/A _11194_/B vssd1 vssd1 vccd1 vccd1 _11194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10145_ _10219_/A1 _18163_/Q _18809_/Q _10215_/S vssd1 vssd1 vccd1 vccd1 _10145_/X
+ sky130_fd_sc_hd__a22o_1
X_17810_ _19490_/CLK _17810_/D vssd1 vssd1 vccd1 vccd1 _17810_/Q sky130_fd_sc_hd__dfxtp_4
X_18790_ _19206_/CLK _18790_/D vssd1 vssd1 vccd1 vccd1 _18790_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17741_ _18641_/Q vssd1 vssd1 vccd1 vccd1 _18641_/D sky130_fd_sc_hd__clkbuf_2
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14953_ _14973_/A1 _13788_/Y _14973_/B1 _18652_/Q _14741_/B vssd1 vssd1 vccd1 vccd1
+ _14953_/X sky130_fd_sc_hd__a221o_1
X_10076_ _11745_/B _10076_/B vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__or2_4
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ _13904_/A _13904_/B vssd1 vssd1 vccd1 vccd1 _13904_/Y sky130_fd_sc_hd__nor2_1
X_17672_ _17672_/A0 _19599_/Q _17689_/S vssd1 vssd1 vccd1 vccd1 _19599_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14884_ _14854_/X _14883_/X _14726_/X vssd1 vssd1 vccd1 vccd1 _14884_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19411_ _19519_/CLK _19411_/D vssd1 vssd1 vccd1 vccd1 _19411_/Q sky130_fd_sc_hd__dfxtp_1
X_16623_ _17723_/A0 _19226_/Q _16623_/S vssd1 vssd1 vccd1 vccd1 _19226_/D sky130_fd_sc_hd__mux2_1
XFILLER_262_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13835_ _13323_/B _13817_/X _13834_/X _13968_/A1 vssd1 vssd1 vccd1 vccd1 _13835_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16554_ _10239_/B _19159_/Q _16554_/S vssd1 vssd1 vccd1 vccd1 _19159_/D sky130_fd_sc_hd__mux2_1
X_19342_ _19470_/CLK _19342_/D vssd1 vssd1 vccd1 vccd1 _19342_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13766_ _13763_/A _12837_/B _13962_/B _11545_/A _13765_/Y vssd1 vssd1 vccd1 vccd1
+ _13766_/X sky130_fd_sc_hd__o221a_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ _10963_/Y _10976_/X _10977_/X vssd1 vssd1 vccd1 vccd1 _10978_/X sky130_fd_sc_hd__o21a_2
X_15505_ _15506_/A _15506_/B vssd1 vssd1 vccd1 vccd1 _15532_/A sky130_fd_sc_hd__nor2_1
X_19273_ _19273_/CLK _19273_/D vssd1 vssd1 vccd1 vccd1 _19273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ _12713_/X _12716_/X _12935_/S vssd1 vssd1 vccd1 vccd1 _12717_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16485_ _17684_/A0 _19092_/Q _16485_/S vssd1 vssd1 vccd1 vccd1 _19092_/D sky130_fd_sc_hd__mux2_1
XFILLER_241_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13697_ _13697_/A _13697_/B vssd1 vssd1 vccd1 vccd1 _14151_/A sky130_fd_sc_hd__xnor2_4
X_18224_ _19618_/CLK _18224_/D vssd1 vssd1 vccd1 vccd1 _18224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15436_ _15456_/D _15436_/B vssd1 vssd1 vccd1 vccd1 _15436_/X sky130_fd_sc_hd__xor2_1
XFILLER_176_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12648_ _10453_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _12648_/X sky130_fd_sc_hd__and2b_1
XFILLER_169_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18155_ _19025_/CLK _18155_/D vssd1 vssd1 vccd1 vccd1 _18155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15367_ _15456_/A _15368_/B vssd1 vssd1 vccd1 vccd1 _15385_/B sky130_fd_sc_hd__or2_1
X_12579_ _12579_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _12579_/Y sky130_fd_sc_hd__nor2_8
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17106_ _17199_/B _17116_/A2 _17105_/X _17106_/C1 vssd1 vssd1 vccd1 vccd1 _19386_/D
+ sky130_fd_sc_hd__o211a_1
X_14318_ _18175_/Q _16602_/A0 _14335_/S vssd1 vssd1 vccd1 vccd1 _18175_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18086_ _18700_/CLK _18086_/D vssd1 vssd1 vccd1 vccd1 _18086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15298_ _15275_/Y _15280_/B _15277_/B vssd1 vssd1 vccd1 vccd1 _15299_/B sky130_fd_sc_hd__o21ai_4
XFILLER_183_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17037_ _19355_/Q _17041_/B vssd1 vssd1 vccd1 vccd1 _17037_/X sky130_fd_sc_hd__or2_1
X_14249_ _18296_/Q _14261_/A2 _14248_/X _14451_/B vssd1 vssd1 vccd1 vccd1 _18122_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout808 _15801_/Y vssd1 vssd1 vccd1 vccd1 _15817_/S sky130_fd_sc_hd__buf_12
XFILLER_140_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout819 _14325_/S vssd1 vssd1 vccd1 vccd1 _14338_/S sky130_fd_sc_hd__buf_8
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _10036_/S _09786_/X _09787_/X vssd1 vssd1 vccd1 vccd1 _09790_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_280_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _19118_/CLK _18988_/D vssd1 vssd1 vccd1 vccd1 _18988_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _18660_/CLK _17939_/D vssd1 vssd1 vccd1 vccd1 _17939_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1390 _09092_/Y vssd1 vssd1 vccd1 vccd1 _09843_/S sky130_fd_sc_hd__buf_8
XFILLER_27_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19609_ _19609_/CLK _19609_/D vssd1 vssd1 vccd1 vccd1 _19609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ _11417_/B1 _09222_/X _09223_/X _09209_/X vssd1 vssd1 vccd1 vccd1 _09224_/X
+ sky130_fd_sc_hd__o31a_4
XFILLER_158_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09155_ _18383_/Q _09908_/B1 _09154_/Y _09992_/A vssd1 vssd1 vccd1 vccd1 _09156_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_163_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09086_ _09086_/A _12023_/A vssd1 vssd1 vccd1 vccd1 _09086_/Y sky130_fd_sc_hd__nor2_8
XFILLER_238_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09988_ _09031_/S _09331_/Y _09987_/Y _09985_/Y vssd1 vssd1 vccd1 vccd1 _09988_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08939_ _08939_/A _08939_/B _08939_/C vssd1 vssd1 vccd1 vccd1 _08947_/A sky130_fd_sc_hd__and3_4
XFILLER_264_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11950_ _11953_/B2 _11904_/B _11953_/A2 input238/X vssd1 vssd1 vccd1 vccd1 _11950_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_229_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _11131_/A _10901_/B _10901_/C vssd1 vssd1 vccd1 vccd1 _10901_/X sky130_fd_sc_hd__or3_1
XFILLER_205_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11881_ _11807_/Y _11875_/Y _11880_/X vssd1 vssd1 vccd1 vccd1 _11882_/C sky130_fd_sc_hd__o21ai_2
XFILLER_264_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13620_ _12732_/S _13229_/X _13232_/Y _13863_/B2 vssd1 vssd1 vccd1 vccd1 _13620_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10832_ _10832_/A _12640_/B vssd1 vssd1 vccd1 vccd1 _11537_/B sky130_fd_sc_hd__and2_4
XFILLER_199_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13551_ _17842_/Q _13846_/B vssd1 vssd1 vccd1 vccd1 _13551_/Y sky130_fd_sc_hd__nor2_1
X_10763_ _10761_/X _10762_/X _11577_/S vssd1 vssd1 vccd1 vccd1 _10763_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ _12502_/A _12554_/B vssd1 vssd1 vccd1 vccd1 _12563_/A sky130_fd_sc_hd__or2_1
XFILLER_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16270_ _17668_/A0 _18884_/Q _16288_/S vssd1 vssd1 vccd1 vccd1 _18884_/D sky130_fd_sc_hd__mux2_1
X_13482_ _13482_/A vssd1 vssd1 vccd1 vccd1 _13482_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ _11173_/S _18801_/Q _11249_/S vssd1 vssd1 vccd1 vccd1 _10694_/X sky130_fd_sc_hd__and3_1
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15221_ _15200_/B _15201_/X _15198_/X vssd1 vssd1 vccd1 vccd1 _15222_/B sky130_fd_sc_hd__o21ai_2
X_12433_ _17887_/Q _12433_/B _12433_/C vssd1 vssd1 vccd1 vccd1 _12433_/X sky130_fd_sc_hd__or3_1
XFILLER_185_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ _15259_/B _12927_/Y _15285_/A3 _15151_/Y vssd1 vssd1 vccd1 vccd1 _15152_/X
+ sky130_fd_sc_hd__a31o_1
X_12364_ _12408_/B _12364_/B vssd1 vssd1 vccd1 vccd1 _12364_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14103_ _16553_/A0 _18043_/Q _14106_/S vssd1 vssd1 vccd1 vccd1 _18043_/D sky130_fd_sc_hd__mux2_1
X_11315_ _19632_/Q _18921_/Q _11325_/S vssd1 vssd1 vccd1 vccd1 _11315_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15083_ _15083_/A _15083_/B vssd1 vssd1 vccd1 vccd1 _15083_/Y sky130_fd_sc_hd__nor2_2
X_12295_ _14680_/B _14672_/C vssd1 vssd1 vccd1 vccd1 _14675_/A sky130_fd_sc_hd__or2_1
XFILLER_154_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14034_ _17982_/Q _14034_/B vssd1 vssd1 vccd1 vccd1 _14034_/X sky130_fd_sc_hd__or2_1
X_18911_ _19622_/CLK _18911_/D vssd1 vssd1 vccd1 vccd1 _18911_/Q sky130_fd_sc_hd__dfxtp_1
X_11246_ _18251_/Q _18826_/Q _11247_/S vssd1 vssd1 vccd1 vccd1 _11246_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18842_ _19639_/CLK _18842_/D vssd1 vssd1 vccd1 vccd1 _18842_/Q sky130_fd_sc_hd__dfxtp_1
X_11177_ _09137_/S _11166_/X _11174_/X _11176_/X vssd1 vssd1 vccd1 vccd1 _11177_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10128_ _18656_/Q _10128_/B vssd1 vssd1 vccd1 vccd1 _10128_/X sky130_fd_sc_hd__or2_1
XFILLER_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15985_ _18708_/Q _16019_/A2 _15984_/X _14197_/A vssd1 vssd1 vccd1 vccd1 _18708_/D
+ sky130_fd_sc_hd__o211a_1
X_18773_ _18775_/CLK _18773_/D vssd1 vssd1 vccd1 vccd1 _18773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14936_ _15006_/A1 _14935_/X _15006_/B1 vssd1 vssd1 vccd1 vccd1 _14936_/Y sky130_fd_sc_hd__o21ai_2
X_17724_ _17724_/A _17724_/B vssd1 vssd1 vccd1 vccd1 _17724_/Y sky130_fd_sc_hd__nor2_1
X_10059_ _11622_/C1 _10053_/X _10056_/X _10058_/X vssd1 vssd1 vccd1 vccd1 _10059_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_250_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18632_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17655_ _17688_/A0 _19583_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _19583_/D sky130_fd_sc_hd__mux2_1
X_14867_ _14867_/A vssd1 vssd1 vccd1 vccd1 _14867_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_250_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16606_ _16606_/A0 _19209_/Q _16618_/S vssd1 vssd1 vccd1 vccd1 _19209_/D sky130_fd_sc_hd__mux2_1
X_13818_ _13818_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13818_/X sky130_fd_sc_hd__or2_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17586_ _19535_/Q _17561_/B _17588_/B1 _17585_/X vssd1 vssd1 vccd1 vccd1 _19535_/D
+ sky130_fd_sc_hd__o211a_1
X_14798_ _18481_/Q _14889_/B1 _14797_/Y _12249_/A vssd1 vssd1 vccd1 vccd1 _18481_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16537_ _17670_/A0 _19142_/Q _16556_/S vssd1 vssd1 vccd1 vccd1 _19142_/D sky130_fd_sc_hd__mux2_1
X_19325_ _19327_/CLK _19325_/D vssd1 vssd1 vccd1 vccd1 _19325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_259_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13749_ _19515_/Q _13947_/A2 _13947_/B1 _13748_/X vssd1 vssd1 vccd1 vccd1 _13749_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16468_ _16501_/A0 _19075_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _19075_/D sky130_fd_sc_hd__mux2_1
X_19256_ _19261_/CLK _19256_/D vssd1 vssd1 vccd1 vccd1 _19256_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_188_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18207_ _19114_/CLK _18207_/D vssd1 vssd1 vccd1 vccd1 _18207_/Q sky130_fd_sc_hd__dfxtp_1
X_15419_ _15419_/A _15419_/B vssd1 vssd1 vccd1 vccd1 _15421_/A sky130_fd_sc_hd__nand2_1
X_19187_ _19219_/CLK _19187_/D vssd1 vssd1 vccd1 vccd1 _19187_/Q sky130_fd_sc_hd__dfxtp_1
X_16399_ _17697_/A0 _19008_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _19008_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18138_ _19608_/CLK _18138_/D vssd1 vssd1 vccd1 vccd1 _18138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18069_ _19226_/CLK _18069_/D vssd1 vssd1 vccd1 vccd1 _18069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09911_ _08946_/B _09904_/Y _09910_/Y _17921_/Q vssd1 vssd1 vccd1 vccd1 _09911_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_160_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout605 _17475_/A2 vssd1 vssd1 vccd1 vccd1 _17445_/A2 sky130_fd_sc_hd__buf_2
Xfanout616 _17558_/B vssd1 vssd1 vccd1 vccd1 _17561_/B sky130_fd_sc_hd__buf_6
Xfanout627 _16947_/S vssd1 vssd1 vccd1 vccd1 _16927_/S sky130_fd_sc_hd__clkbuf_4
X_09842_ _18628_/Q _18050_/Q _11160_/S vssd1 vssd1 vccd1 vccd1 _09842_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout638 _17337_/S vssd1 vssd1 vccd1 vccd1 _17379_/S sky130_fd_sc_hd__buf_8
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout649 _17073_/B vssd1 vssd1 vccd1 vccd1 _17077_/B sky130_fd_sc_hd__buf_2
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09773_ _09086_/A _09750_/X _09772_/X _09107_/D vssd1 vssd1 vccd1 vccd1 _09773_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_273_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09207_ _09205_/X _09206_/X _10225_/S vssd1 vssd1 vccd1 vccd1 _09207_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09138_ _09116_/X _09124_/X _09137_/X _10260_/B1 vssd1 vssd1 vccd1 vccd1 _09138_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_120_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09069_ _09083_/A vssd1 vssd1 vccd1 vccd1 _11706_/C sky130_fd_sc_hd__inv_8
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11100_ _09107_/D _11089_/X _11097_/X _11099_/X vssd1 vssd1 vccd1 vccd1 _11100_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_265_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12080_ _17915_/Q _12088_/A2 _12079_/X _17419_/C1 vssd1 vssd1 vccd1 vccd1 _17817_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11031_ _11029_/X _11030_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _11031_/X sky130_fd_sc_hd__mux2_1
XFILLER_249_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15770_ _15770_/A _15770_/B vssd1 vssd1 vccd1 vccd1 _15770_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_40_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12982_ _15330_/A _12982_/B vssd1 vssd1 vccd1 vccd1 _12982_/Y sky130_fd_sc_hd__nor2_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _18473_/Q _14720_/A _14720_/Y _17330_/A vssd1 vssd1 vccd1 vccd1 _18473_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11933_ _11953_/B2 _11827_/B _11827_/C _11953_/A2 input219/X vssd1 vssd1 vccd1 vccd1
+ _11933_/X sky130_fd_sc_hd__a32o_4
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_510 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_521 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_532 _18396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _13224_/A _15118_/A _17445_/B1 _17800_/Q _17445_/C1 vssd1 vssd1 vccd1 vccd1
+ _17440_/X sky130_fd_sc_hd__a221o_1
XFILLER_261_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _17711_/A0 _18458_/Q _14664_/S vssd1 vssd1 vccd1 vccd1 _18458_/D sky130_fd_sc_hd__mux2_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11864_ _11864_/A _11864_/B vssd1 vssd1 vccd1 vccd1 _11901_/A sky130_fd_sc_hd__or2_2
XANTENNA_543 _18109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13603_ _13966_/C1 _13601_/X _13602_/X _13599_/Y vssd1 vssd1 vccd1 vccd1 _13603_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _18864_/Q _10815_/B vssd1 vssd1 vccd1 vccd1 _10815_/X sky130_fd_sc_hd__or2_1
X_17371_ _19483_/Q _17202_/B _17379_/S vssd1 vssd1 vccd1 vccd1 _17372_/B sky130_fd_sc_hd__mux2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _18400_/Q _14589_/A2 _14589_/B1 input29/X vssd1 vssd1 vccd1 vccd1 _14584_/B
+ sky130_fd_sc_hd__o22a_1
X_11795_ _11799_/A _11799_/B _11820_/B vssd1 vssd1 vccd1 vccd1 _11795_/X sky130_fd_sc_hd__and3_1
XFILLER_198_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19110_ _19142_/CLK _19110_/D vssd1 vssd1 vccd1 vccd1 _19110_/Q sky130_fd_sc_hd__dfxtp_1
X_16322_ _17720_/A0 _18935_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _18935_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13534_ _13958_/B _14147_/B _13892_/B1 vssd1 vssd1 vccd1 vccd1 _13534_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_201_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10746_ _10742_/X _10745_/X _10746_/S vssd1 vssd1 vccd1 vccd1 _10746_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19041_ _19624_/CLK _19041_/D vssd1 vssd1 vccd1 vccd1 _19041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16253_ _17717_/A0 _18868_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _18868_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_147_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19552_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_201_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13465_ _13465_/A _13465_/B _13465_/C vssd1 vssd1 vccd1 vccd1 _13466_/B sky130_fd_sc_hd__and3_1
XFILLER_145_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ _10677_/A _12729_/A vssd1 vssd1 vccd1 vccd1 _11541_/B sky130_fd_sc_hd__and2_4
X_15204_ _15204_/A _15204_/B vssd1 vssd1 vccd1 vccd1 _15204_/Y sky130_fd_sc_hd__xnor2_1
X_12416_ _17913_/Q _12427_/A _12415_/Y _12428_/C1 vssd1 vssd1 vccd1 vccd1 _17913_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16184_ _17714_/A0 _18801_/Q _16189_/S vssd1 vssd1 vccd1 vccd1 _18801_/D sky130_fd_sc_hd__mux2_1
X_13396_ _13323_/X _13384_/X _13395_/X _13968_/B2 vssd1 vssd1 vccd1 vccd1 _13396_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15135_ _15135_/A _15135_/B vssd1 vssd1 vccd1 vccd1 _15137_/B sky130_fd_sc_hd__xor2_2
X_12347_ _17890_/Q _12349_/A _12346_/Y _12350_/C1 vssd1 vssd1 vccd1 vccd1 _17890_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15066_ _18550_/Q _17677_/A0 _15078_/S vssd1 vssd1 vccd1 vccd1 _18550_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12278_ _18091_/Q _12305_/A2 _12305_/B1 _18514_/Q vssd1 vssd1 vccd1 vccd1 _12474_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14017_ _17973_/Q _14020_/B _14016_/Y _14037_/C1 vssd1 vssd1 vccd1 vccd1 _17973_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11229_ _11250_/A1 _19146_/Q _11226_/S _19114_/Q _11567_/S vssd1 vssd1 vccd1 vccd1
+ _11229_/X sky130_fd_sc_hd__o221a_1
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18825_ _19632_/CLK _18825_/D vssd1 vssd1 vccd1 vccd1 _18825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18756_ _18775_/CLK _18756_/D vssd1 vssd1 vccd1 vccd1 _18756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15968_ _18699_/Q _15970_/A2 _15976_/B1 _18748_/Q _15976_/C1 vssd1 vssd1 vccd1 vccd1
+ _15968_/X sky130_fd_sc_hd__a221o_1
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17707_ _17707_/A0 _19633_/Q _17718_/S vssd1 vssd1 vccd1 vccd1 _19633_/D sky130_fd_sc_hd__mux2_1
XFILLER_264_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14919_ _14915_/Y _14918_/X _14950_/B1 vssd1 vssd1 vccd1 vccd1 _14919_/Y sky130_fd_sc_hd__a21oi_4
X_15899_ _15899_/A _15941_/S _15905_/C vssd1 vssd1 vccd1 vccd1 _15899_/X sky130_fd_sc_hd__and3_1
X_18687_ _19276_/CLK _18687_/D vssd1 vssd1 vccd1 vccd1 _18687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17638_ _17671_/A0 _19566_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _19566_/D sky130_fd_sc_hd__mux2_1
XFILLER_247_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17569_ _17569_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17569_/X sky130_fd_sc_hd__or2_1
X_19308_ _19310_/CLK _19308_/D vssd1 vssd1 vccd1 vccd1 _19308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19239_ _19273_/CLK _19239_/D vssd1 vssd1 vccd1 vccd1 _19239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09825_ _17954_/Q _11216_/A2 _08947_/X _17922_/Q _09824_/X vssd1 vssd1 vccd1 vccd1
+ _09825_/X sky130_fd_sc_hd__a221o_4
XFILLER_247_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09756_ _11565_/A1 _19557_/Q _09770_/S _19589_/Q vssd1 vssd1 vccd1 vccd1 _09756_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_274_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09687_ _18443_/Q _18344_/Q _09688_/S vssd1 vssd1 vccd1 vccd1 _09687_/X sky130_fd_sc_hd__mux2_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ _18125_/Q _10599_/Y _13739_/A vssd1 vssd1 vccd1 vccd1 _12650_/B sky130_fd_sc_hd__mux2_4
X_11580_ _11584_/A1 _19226_/Q _19194_/Q _11581_/S _09095_/A vssd1 vssd1 vccd1 vccd1
+ _11580_/X sky130_fd_sc_hd__a221o_1
XFILLER_80_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ _17944_/Q _11451_/A2 _10530_/X vssd1 vssd1 vccd1 vccd1 _10531_/X sky130_fd_sc_hd__o21a_4
XFILLER_183_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ _17833_/Q _13944_/B _13248_/X _13249_/X vssd1 vssd1 vccd1 vccd1 _13250_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10462_ _10460_/X _10461_/X _10633_/A vssd1 vssd1 vccd1 vccd1 _10462_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12201_ _12203_/A _12201_/B _12202_/B vssd1 vssd1 vccd1 vccd1 _17864_/D sky130_fd_sc_hd__nor3_1
XFILLER_182_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13181_ _13167_/A _12768_/A _12583_/Y vssd1 vssd1 vccd1 vccd1 _13181_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10393_ _18620_/Q _18191_/Q _11576_/S vssd1 vssd1 vccd1 vccd1 _10393_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12132_ _17838_/Q _12130_/B _12131_/Y vssd1 vssd1 vccd1 vccd1 _17838_/D sky130_fd_sc_hd__o21a_1
XFILLER_2_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16940_ _17346_/A _16940_/B vssd1 vssd1 vccd1 vccd1 _19319_/D sky130_fd_sc_hd__and2_1
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12063_ _17809_/Q _12085_/B vssd1 vssd1 vccd1 vccd1 _12063_/X sky130_fd_sc_hd__or2_1
Xfanout1901 _14991_/C1 vssd1 vssd1 vccd1 vccd1 _16740_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_284_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11014_ _11469_/A1 _18612_/Q _18183_/Q _11477_/S vssd1 vssd1 vccd1 vccd1 _11014_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16871_ _19302_/Q _17571_/A _16927_/S vssd1 vssd1 vccd1 vccd1 _16872_/B sky130_fd_sc_hd__mux2_1
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout980 _13427_/A1 vssd1 vssd1 vccd1 vccd1 _13303_/B2 sky130_fd_sc_hd__buf_6
XFILLER_237_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18610_ _19634_/CLK _18610_/D vssd1 vssd1 vccd1 vccd1 _18610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _18614_/Q _16314_/A0 _15833_/S vssd1 vssd1 vccd1 vccd1 _18614_/D sky130_fd_sc_hd__mux2_1
Xfanout991 _11647_/X vssd1 vssd1 vccd1 vccd1 _11845_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ _19592_/CLK _19590_/D vssd1 vssd1 vccd1 vccd1 _19590_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18541_ _19595_/CLK _18541_/D vssd1 vssd1 vccd1 vccd1 _18541_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _19485_/Q _19419_/Q vssd1 vssd1 vccd1 vccd1 _15753_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12965_ _19236_/Q _13495_/A2 _13495_/B1 _19268_/Q vssd1 vssd1 vccd1 vccd1 _12965_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ _18570_/Q _11918_/A2 _11706_/B _13147_/A vssd1 vssd1 vccd1 vccd1 _11916_/X
+ sky130_fd_sc_hd__a22o_4
X_14704_ _18102_/Q _14893_/S vssd1 vssd1 vccd1 vccd1 _14704_/X sky130_fd_sc_hd__or2_1
X_18472_ _19229_/CLK _18472_/D vssd1 vssd1 vccd1 vccd1 _18472_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15684_ _15684_/A _15684_/B vssd1 vssd1 vccd1 vccd1 _15685_/A sky130_fd_sc_hd__or2_1
XFILLER_46_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _13046_/A1 _12895_/Y _12745_/X vssd1 vssd1 vccd1 vccd1 _12896_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_340 _11482_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_351 _09854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _17423_/A _17423_/B vssd1 vssd1 vccd1 vccd1 _17423_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_362 _10471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _17661_/A0 _18441_/Q _14648_/S vssd1 vssd1 vccd1 vccd1 _18441_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ _11824_/A _11812_/X _11846_/Y _11826_/A vssd1 vssd1 vccd1 vccd1 _11847_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_373 _18274_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_384 _17587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_395 _09108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _17354_/A _17354_/B vssd1 vssd1 vccd1 vccd1 _19474_/D sky130_fd_sc_hd__and2_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _14576_/A _14566_/B vssd1 vssd1 vccd1 vccd1 _18391_/D sky130_fd_sc_hd__or2_1
X_11778_ _15039_/B _11777_/Y _11726_/B vssd1 vssd1 vccd1 vccd1 _11778_/X sky130_fd_sc_hd__a21o_1
XFILLER_202_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16305_ _17670_/A0 _18918_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _18918_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13517_ _17841_/Q _13846_/B _12548_/X vssd1 vssd1 vccd1 vccd1 _13517_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10729_ _10719_/S _10721_/X _10720_/X _11198_/S vssd1 vssd1 vccd1 vccd1 _10729_/X
+ sky130_fd_sc_hd__a211o_1
X_17285_ _17285_/A _17285_/B vssd1 vssd1 vccd1 vccd1 _19445_/D sky130_fd_sc_hd__nor2_1
X_14497_ _17699_/A0 _18347_/Q _14517_/S vssd1 vssd1 vccd1 vccd1 _18347_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16236_ _17700_/A0 _18851_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _18851_/D sky130_fd_sc_hd__mux2_1
X_19024_ _19607_/CLK _19024_/D vssd1 vssd1 vccd1 vccd1 _19024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13448_ _19248_/Q _13495_/A2 _13495_/B1 _19280_/Q vssd1 vssd1 vccd1 vccd1 _13448_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_162_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16167_ _16597_/A0 _18784_/Q _16189_/S vssd1 vssd1 vccd1 vccd1 _18784_/D sky130_fd_sc_hd__mux2_1
X_13379_ _17869_/Q _13847_/A2 _13854_/B1 _13378_/X vssd1 vssd1 vccd1 vccd1 _13379_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15118_ _15118_/A _15118_/B vssd1 vssd1 vccd1 vccd1 _15118_/Y sky130_fd_sc_hd__nand2_1
X_16098_ _16142_/A1 _16097_/Y _16149_/A vssd1 vssd1 vccd1 vccd1 _18751_/D sky130_fd_sc_hd__a21oi_1
XFILLER_173_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15049_ _18533_/Q _17660_/A0 _15076_/S vssd1 vssd1 vccd1 vccd1 _18533_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19623_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_205_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09610_ _09948_/B _15194_/A _09562_/X vssd1 vssd1 vccd1 vccd1 _12614_/B sky130_fd_sc_hd__a21boi_4
X_18808_ _19647_/CLK _18808_/D vssd1 vssd1 vccd1 vccd1 _18808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09541_ _18242_/Q _18817_/Q _09542_/S vssd1 vssd1 vccd1 vccd1 _09541_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18739_ _18741_/CLK _18739_/D vssd1 vssd1 vccd1 vccd1 _18739_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09472_ _11257_/C1 _11800_/C _11800_/D _11411_/A vssd1 vssd1 vccd1 vccd1 _09472_/X
+ sky130_fd_sc_hd__a31o_1
XPHY_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1208 _12667_/X vssd1 vssd1 vccd1 vccd1 _12712_/S sky130_fd_sc_hd__buf_2
XFILLER_266_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1219 _12448_/C vssd1 vssd1 vccd1 vccd1 _13971_/A2 sky130_fd_sc_hd__buf_6
XFILLER_59_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09808_ _11282_/A _09806_/X _09807_/X _11285_/S vssd1 vssd1 vccd1 vccd1 _09808_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_15__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09739_ _11691_/B1 _09907_/A _09738_/X _11692_/A1 _18376_/Q vssd1 vssd1 vccd1 vccd1
+ _09739_/X sky130_fd_sc_hd__o32a_1
XFILLER_216_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12750_ _12936_/S _12749_/X _12746_/X vssd1 vssd1 vccd1 vccd1 _12750_/X sky130_fd_sc_hd__o21a_1
XFILLER_216_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _14346_/B _11701_/B _11701_/C _11701_/D vssd1 vssd1 vccd1 vccd1 _11701_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12681_ _12594_/B _12597_/B _12835_/A vssd1 vssd1 vccd1 vccd1 _12681_/X sky130_fd_sc_hd__mux2_4
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _19229_/Q _15014_/B _18274_/D vssd1 vssd1 vccd1 vccd1 _18271_/D sky130_fd_sc_hd__and3_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _13938_/B _13958_/A vssd1 vssd1 vccd1 vccd1 _11728_/A sky130_fd_sc_hd__and2_1
XFILLER_168_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ _14351_/A _16459_/C vssd1 vssd1 vccd1 vccd1 _14351_/Y sky130_fd_sc_hd__nor2_8
XFILLER_211_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11563_ _11568_/A _11562_/X _11563_/B1 vssd1 vssd1 vccd1 vccd1 _11563_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13302_ _19372_/Q _13301_/X _13925_/S vssd1 vssd1 vccd1 vccd1 _13302_/X sky130_fd_sc_hd__mux2_2
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17070_ _17575_/A _17114_/A2 _17069_/X _17559_/A vssd1 vssd1 vccd1 vccd1 _19368_/D
+ sky130_fd_sc_hd__o211a_1
X_10514_ _10510_/X _10513_/X _12320_/B vssd1 vssd1 vccd1 vccd1 _10514_/X sky130_fd_sc_hd__mux2_1
X_14282_ _16203_/A0 _18141_/Q _14301_/S vssd1 vssd1 vccd1 vccd1 _18141_/D sky130_fd_sc_hd__mux2_1
X_11494_ _11492_/X _11493_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _11494_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16021_ _16020_/A _16056_/B _18726_/Q vssd1 vssd1 vccd1 vccd1 _16021_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13233_ _13863_/B2 _13229_/X _13232_/Y _12712_/S vssd1 vssd1 vccd1 vccd1 _13233_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ _10663_/S _10432_/X _10433_/X vssd1 vssd1 vccd1 vccd1 _10445_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164_ _17831_/Q _13164_/A2 _13164_/B1 _17863_/Q vssd1 vssd1 vccd1 vccd1 _13164_/X
+ sky130_fd_sc_hd__a22o_1
X_10376_ _11210_/A1 _10341_/A2 _10375_/Y _11055_/B2 vssd1 vssd1 vccd1 vccd1 _13818_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12115_ _12203_/A _12120_/C vssd1 vssd1 vccd1 vccd1 _12115_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17972_ _18700_/CLK _17972_/D vssd1 vssd1 vccd1 vccd1 _17972_/Q sky130_fd_sc_hd__dfxtp_1
X_13095_ _09560_/X _13316_/B _12836_/Y _13083_/A _13260_/A vssd1 vssd1 vccd1 vccd1
+ _13095_/Y sky130_fd_sc_hd__a221oi_4
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16923_ _19315_/Q _17178_/B _16927_/S vssd1 vssd1 vccd1 vccd1 _16924_/B sky130_fd_sc_hd__mux2_1
X_12046_ _17898_/Q _12052_/A2 _12045_/X _13100_/A vssd1 vssd1 vccd1 vccd1 _17800_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1720 _18739_/Q vssd1 vssd1 vccd1 vccd1 _16054_/A sky130_fd_sc_hd__buf_4
Xfanout1731 _15088_/B vssd1 vssd1 vccd1 vccd1 _15086_/B sky130_fd_sc_hd__buf_4
XFILLER_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1742 _18273_/Q vssd1 vssd1 vccd1 vccd1 _14844_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1753 _11583_/A vssd1 vssd1 vccd1 vccd1 _11328_/S sky130_fd_sc_hd__buf_8
XFILLER_78_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1764 _15129_/B2 vssd1 vssd1 vccd1 vccd1 _12320_/A sky130_fd_sc_hd__buf_12
X_19642_ _19642_/CLK _19642_/D vssd1 vssd1 vccd1 vccd1 _19642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1775 _17909_/Q vssd1 vssd1 vccd1 vccd1 _12471_/A0 sky130_fd_sc_hd__buf_12
X_16854_ _19298_/Q _17563_/A _16967_/S vssd1 vssd1 vccd1 vccd1 _16855_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1786 _17905_/Q vssd1 vssd1 vccd1 vccd1 _08896_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1797 _08816_/A vssd1 vssd1 vccd1 vccd1 _08991_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15805_ _18597_/Q _16595_/A0 _15817_/S vssd1 vssd1 vccd1 vccd1 _18597_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19573_ _19573_/CLK _19573_/D vssd1 vssd1 vccd1 vccd1 _19573_/Q sky130_fd_sc_hd__dfxtp_1
X_16785_ _19283_/Q _16786_/B vssd1 vssd1 vccd1 vccd1 _16787_/B sky130_fd_sc_hd__nor2_1
X_13997_ _17963_/Q _14032_/B _13996_/Y _16153_/D vssd1 vssd1 vccd1 vccd1 _17963_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18524_ _19286_/CLK _18524_/D vssd1 vssd1 vccd1 vccd1 _18524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15736_ _15757_/A _15756_/A vssd1 vssd1 vccd1 vccd1 _15738_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12948_ _11734_/B _14155_/B _13358_/A1 vssd1 vssd1 vccd1 vccd1 _12948_/X sky130_fd_sc_hd__o21a_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_162_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19540_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18455_ _19634_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_170 _13213_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ _13039_/S _12879_/B vssd1 vssd1 vccd1 vccd1 _12879_/Y sky130_fd_sc_hd__nor2_1
X_15667_ _15690_/A _15664_/Y _15666_/Y _15751_/A vssd1 vssd1 vccd1 vccd1 _15667_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _13546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_192 _14026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17406_ _12956_/A _15118_/A _15117_/A _17793_/Q _15116_/B vssd1 vssd1 vccd1 vccd1
+ _17406_/X sky130_fd_sc_hd__a221o_1
X_14618_ _17677_/A0 _18425_/Q _14630_/S vssd1 vssd1 vccd1 vccd1 _18425_/D sky130_fd_sc_hd__mux2_1
XFILLER_194_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15598_ _15787_/A _15639_/B vssd1 vssd1 vccd1 vccd1 _15638_/C sky130_fd_sc_hd__xnor2_4
X_18386_ _19471_/CLK _18386_/D vssd1 vssd1 vccd1 vccd1 _18386_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14549_ _18383_/Q _14575_/A2 _14575_/B1 input11/X vssd1 vssd1 vccd1 vccd1 _14550_/B
+ sky130_fd_sc_hd__o22a_1
X_17337_ _19466_/Q _17579_/A _17337_/S vssd1 vssd1 vccd1 vccd1 _17338_/B sky130_fd_sc_hd__mux2_1
XFILLER_187_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17268_ _19440_/Q _17313_/B vssd1 vssd1 vccd1 vccd1 _17268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19007_ _19138_/CLK _19007_/D vssd1 vssd1 vccd1 vccd1 _19007_/Q sky130_fd_sc_hd__dfxtp_1
X_16219_ _17716_/A0 _18835_/Q _16226_/S vssd1 vssd1 vccd1 vccd1 _18835_/D sky130_fd_sc_hd__mux2_1
X_17199_ _17199_/A _17199_/B vssd1 vssd1 vccd1 vccd1 _17199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08972_ _10419_/S _08972_/B vssd1 vssd1 vccd1 vccd1 _08977_/A sky130_fd_sc_hd__and2_1
XFILLER_142_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09524_ _11210_/A1 _15808_/A1 _09523_/X vssd1 vssd1 vccd1 vccd1 _15214_/A sky130_fd_sc_hd__a21oi_4
XFILLER_25_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09455_ _19042_/Q _19010_/Q _09464_/S vssd1 vssd1 vccd1 vccd1 _09455_/X sky130_fd_sc_hd__mux2_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09386_ _09384_/X _09385_/X _10200_/S vssd1 vssd1 vccd1 vccd1 _09386_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10230_ _18130_/Q _13874_/A _13904_/A vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__mux2_4
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10161_ _12656_/A vssd1 vssd1 vccd1 vccd1 _13908_/A sky130_fd_sc_hd__inv_6
XFILLER_133_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput380 _11933_/X vssd1 vssd1 vccd1 vccd1 din0[13] sky130_fd_sc_hd__buf_4
XFILLER_267_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1005 _10081_/X vssd1 vssd1 vccd1 vccd1 _11181_/B1 sky130_fd_sc_hd__buf_6
Xoutput391 _11943_/X vssd1 vssd1 vccd1 vccd1 din0[23] sky130_fd_sc_hd__buf_4
XFILLER_273_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1016 _14412_/S vssd1 vssd1 vccd1 vccd1 _14415_/S sky130_fd_sc_hd__buf_12
XFILLER_0_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1027 _16530_/A0 vssd1 vssd1 vccd1 vccd1 _17696_/A0 sky130_fd_sc_hd__clkbuf_4
X_10092_ _10090_/X _10091_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _10093_/B sky130_fd_sc_hd__mux2_1
Xfanout1038 _09491_/X vssd1 vssd1 vccd1 vccd1 _17698_/A0 sky130_fd_sc_hd__buf_2
XFILLER_48_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1049 _17528_/B vssd1 vssd1 vccd1 vccd1 _17437_/A2 sky130_fd_sc_hd__buf_6
XFILLER_247_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13920_ _17885_/Q _13945_/A2 _13919_/X _13920_/B2 _13952_/B1 vssd1 vssd1 vccd1 vccd1
+ _13920_/X sky130_fd_sc_hd__a221o_1
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13851_ _19452_/Q _13949_/A2 _13849_/X _13850_/X _13949_/C1 vssd1 vssd1 vccd1 vccd1
+ _13851_/X sky130_fd_sc_hd__o221a_1
XFILLER_274_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12802_ _12800_/X _12938_/B _12933_/A vssd1 vssd1 vccd1 vccd1 _12803_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16570_ _09105_/A _19174_/Q _16589_/S vssd1 vssd1 vccd1 vccd1 _19174_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13782_ _19418_/Q _13948_/A2 _13948_/B1 vssd1 vssd1 vccd1 vccd1 _13782_/X sky130_fd_sc_hd__a21o_1
X_10994_ _11469_/A1 _18222_/Q _11386_/S _18957_/Q _11464_/C1 vssd1 vssd1 vccd1 vccd1
+ _10994_/X sky130_fd_sc_hd__o221a_1
XFILLER_203_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12733_ _12599_/B _12640_/B _12733_/S vssd1 vssd1 vccd1 vccd1 _12734_/B sky130_fd_sc_hd__mux2_1
X_15521_ _15519_/Y _15521_/B vssd1 vssd1 vccd1 vccd1 _15522_/B sky130_fd_sc_hd__nand2b_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18240_ _19619_/CLK _18240_/D vssd1 vssd1 vccd1 vccd1 _18240_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _15452_/A _15452_/B vssd1 vssd1 vccd1 vccd1 _15452_/Y sky130_fd_sc_hd__nand2_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12664_ _11629_/B _12663_/B _11627_/Y vssd1 vssd1 vccd1 vccd1 _14155_/A sky130_fd_sc_hd__a21oi_2
XFILLER_230_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _17710_/A0 _18254_/Q _14415_/S vssd1 vssd1 vccd1 vccd1 _18254_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11615_ _19130_/Q _19162_/Q _11617_/S vssd1 vssd1 vccd1 vccd1 _11615_/X sky130_fd_sc_hd__mux2_1
X_18171_ _18632_/CLK _18171_/D vssd1 vssd1 vccd1 vccd1 _18171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15383_ _17901_/Q _15429_/A2 _15484_/A vssd1 vssd1 vccd1 vccd1 _15387_/B sky130_fd_sc_hd__o21a_1
X_12595_ _12595_/A _12595_/B vssd1 vssd1 vccd1 vccd1 _12595_/Y sky130_fd_sc_hd__nor2_2
XFILLER_156_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14334_ _18191_/Q _17718_/A0 _14339_/S vssd1 vssd1 vccd1 vccd1 _18191_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17122_ _19392_/Q _17120_/Y _17121_/X vssd1 vssd1 vccd1 vccd1 _19392_/D sky130_fd_sc_hd__o21ba_1
X_11546_ _12647_/B vssd1 vssd1 vccd1 vccd1 _13763_/A sky130_fd_sc_hd__inv_2
XFILLER_184_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17053_ _19360_/Q _17113_/B vssd1 vssd1 vccd1 vccd1 _17053_/X sky130_fd_sc_hd__or2_1
XFILLER_167_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14265_ _18304_/Q _14267_/A2 _14264_/X _14451_/B vssd1 vssd1 vccd1 vccd1 _18130_/D
+ sky130_fd_sc_hd__o211a_1
X_11477_ _18606_/Q _18177_/Q _11477_/S vssd1 vssd1 vccd1 vccd1 _11477_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16004_ _18717_/Q _16016_/A2 _16004_/B1 _18766_/Q _16004_/C1 vssd1 vssd1 vccd1 vccd1
+ _16004_/X sky130_fd_sc_hd__a221o_1
X_13216_ _17832_/Q _13944_/B _13214_/X _13215_/X vssd1 vssd1 vccd1 vccd1 _13216_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_171_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10428_ _11511_/A _10426_/X _10427_/X _11507_/S vssd1 vssd1 vccd1 vccd1 _10428_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14196_ _18709_/Q _18096_/Q _14200_/S vssd1 vssd1 vccd1 vccd1 _14197_/B sky130_fd_sc_hd__mux2_1
XFILLER_171_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13147_/A _13224_/B vssd1 vssd1 vccd1 vccd1 _13147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10359_ _19062_/Q _19030_/Q _10370_/S vssd1 vssd1 vccd1 vccd1 _10359_/X sky130_fd_sc_hd__mux2_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _17958_/CLK _17955_/D vssd1 vssd1 vccd1 vccd1 _17955_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13078_ _13438_/A _13058_/X _13563_/B1 vssd1 vssd1 vccd1 vccd1 _13079_/C sky130_fd_sc_hd__a21o_1
XFILLER_140_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _16848_/S _17935_/Q _16905_/X vssd1 vssd1 vccd1 vccd1 _17589_/A sky130_fd_sc_hd__o21a_4
Xfanout1550 _10280_/S vssd1 vssd1 vccd1 vccd1 _10300_/S sky130_fd_sc_hd__buf_6
X_12029_ _12029_/A _12035_/B vssd1 vssd1 vccd1 vccd1 _12029_/Y sky130_fd_sc_hd__nand2_1
Xfanout1561 _11286_/B1 vssd1 vssd1 vccd1 vccd1 _11608_/C1 sky130_fd_sc_hd__buf_6
XFILLER_272_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17886_ _19327_/CLK _17886_/D vssd1 vssd1 vccd1 vccd1 _17886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1572 _10653_/C1 vssd1 vssd1 vccd1 vccd1 _11127_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_254_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1583 _10881_/S1 vssd1 vssd1 vccd1 vccd1 _11338_/S1 sky130_fd_sc_hd__buf_4
XFILLER_265_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19625_ _19625_/CLK _19625_/D vssd1 vssd1 vccd1 vccd1 _19625_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1594 _08894_/Y vssd1 vssd1 vccd1 vccd1 _11622_/C1 sky130_fd_sc_hd__clkbuf_8
X_16837_ _16821_/A _17820_/Q _12483_/Y vssd1 vssd1 vccd1 vccd1 _17052_/C sky130_fd_sc_hd__a21o_1
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19556_ _19588_/CLK _19556_/D vssd1 vssd1 vccd1 vccd1 _19556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16768_ _16768_/A _16768_/B _16770_/B vssd1 vssd1 vccd1 vccd1 _19276_/D sky130_fd_sc_hd__nor3_1
XFILLER_222_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18507_ _19229_/CLK _18507_/D vssd1 vssd1 vccd1 vccd1 _18507_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15719_ _13868_/Y _15110_/X _13843_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _15719_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_280_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19487_ _19519_/CLK _19487_/D vssd1 vssd1 vccd1 vccd1 _19487_/Q sky130_fd_sc_hd__dfxtp_2
X_16699_ _19252_/Q _19251_/Q _19250_/Q _16699_/D vssd1 vssd1 vccd1 vccd1 _16708_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_222_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09240_ _09027_/A _10085_/B _09234_/Y _09030_/X vssd1 vssd1 vccd1 vccd1 _09240_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18438_ _19134_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09171_ _11469_/A1 _19564_/Q _09179_/B _19596_/Q _10338_/A1 vssd1 vssd1 vccd1 vccd1
+ _09171_/X sky130_fd_sc_hd__o221a_1
X_18369_ _19648_/CLK _18369_/D vssd1 vssd1 vccd1 vccd1 _18369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput108 dout1[10] vssd1 vssd1 vccd1 vccd1 input108/X sky130_fd_sc_hd__clkbuf_2
X_08955_ _08903_/A _14488_/C _14074_/C _09498_/S _08954_/A vssd1 vssd1 vccd1 vccd1
+ _08956_/D sky130_fd_sc_hd__o221a_1
Xinput119 dout1[20] vssd1 vssd1 vccd1 vccd1 input119/X sky130_fd_sc_hd__clkbuf_2
XFILLER_248_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08886_ _18589_/Q _18588_/Q _18587_/Q _18586_/Q vssd1 vssd1 vccd1 vccd1 _08887_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_257_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09507_ _08896_/A _09506_/X _09501_/X _11515_/B1 vssd1 vssd1 vccd1 vccd1 _09523_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_213_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09438_ _18978_/Q _11167_/B vssd1 vssd1 vccd1 vccd1 _09438_/X sky130_fd_sc_hd__or2_1
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09369_ _10219_/A1 _19203_/Q _19171_/Q _10141_/S _10293_/B1 vssd1 vssd1 vccd1 vccd1
+ _09369_/X sky130_fd_sc_hd__a221o_1
XFILLER_185_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11400_ _18249_/Q _11395_/C _10409_/A _11399_/X vssd1 vssd1 vccd1 vccd1 _11400_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12380_ _17901_/Q _12382_/A _12379_/Y _12383_/C1 vssd1 vssd1 vccd1 vccd1 _17901_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_70 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_81 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _11588_/B1 _11328_/X _11321_/X _09107_/D vssd1 vssd1 vccd1 vccd1 _11331_/X
+ sky130_fd_sc_hd__a211o_2
XANTENNA_92 _10760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14050_ _17667_/A0 _17992_/Q _14072_/S vssd1 vssd1 vccd1 vccd1 _17992_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11262_ _18547_/Q _18422_/Q _18031_/Q _17999_/Q _11284_/B2 _11622_/A1 vssd1 vssd1
+ vccd1 vccd1 _11262_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13001_ _13046_/A1 _12932_/B _12745_/X vssd1 vssd1 vccd1 vccd1 _13001_/Y sky130_fd_sc_hd__o21ai_4
X_10213_ _10219_/A1 _19224_/Q _19192_/Q _10215_/S _10293_/B1 vssd1 vssd1 vccd1 vccd1
+ _10213_/X sky130_fd_sc_hd__a221o_1
XFILLER_134_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11193_ _09723_/S _11192_/X _11508_/B1 vssd1 vssd1 vccd1 vccd1 _11194_/B sky130_fd_sc_hd__a21o_1
XFILLER_134_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10144_ _18873_/Q _10215_/S _10144_/B1 vssd1 vssd1 vccd1 vccd1 _10144_/X sky130_fd_sc_hd__o21a_1
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17740_ _18640_/Q vssd1 vssd1 vccd1 vccd1 _18640_/D sky130_fd_sc_hd__clkbuf_2
X_14952_ _17816_/Q _14982_/B vssd1 vssd1 vccd1 vccd1 _14952_/X sky130_fd_sc_hd__or2_1
X_10075_ _11742_/B _10074_/B _11745_/A vssd1 vssd1 vccd1 vccd1 _10076_/B sky130_fd_sc_hd__a21oi_1
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ _15330_/A _13903_/B vssd1 vssd1 vccd1 vccd1 _13903_/X sky130_fd_sc_hd__or2_1
X_17671_ _17671_/A0 _19598_/Q _17689_/S vssd1 vssd1 vccd1 vccd1 _19598_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14883_ _18120_/Q _14882_/X _14893_/S vssd1 vssd1 vccd1 vccd1 _14883_/X sky130_fd_sc_hd__mux2_2
XFILLER_130_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19410_ _19519_/CLK _19410_/D vssd1 vssd1 vccd1 vccd1 _19410_/Q sky130_fd_sc_hd__dfxtp_2
X_16622_ _16622_/A0 _19225_/Q _16622_/S vssd1 vssd1 vccd1 vccd1 _19225_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13834_ _13931_/A _13832_/X _13833_/Y _13810_/A _13294_/A vssd1 vssd1 vccd1 vccd1
+ _13834_/X sky130_fd_sc_hd__o32a_1
XFILLER_223_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19341_ _19534_/CLK _19341_/D vssd1 vssd1 vccd1 vccd1 _19341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_262_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16553_ _16553_/A0 _19158_/Q _16556_/S vssd1 vssd1 vccd1 vccd1 _19158_/D sky130_fd_sc_hd__mux2_1
X_13765_ _11545_/B _13912_/A2 _14153_/A vssd1 vssd1 vccd1 vccd1 _13765_/Y sky130_fd_sc_hd__a21oi_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10977_ _11131_/A _10977_/B _10977_/C vssd1 vssd1 vccd1 vccd1 _10977_/X sky130_fd_sc_hd__or3_1
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15504_ _18119_/Q _15786_/A2 _15503_/X _15452_/A vssd1 vssd1 vccd1 vccd1 _15506_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_19272_ _19273_/CLK _19272_/D vssd1 vssd1 vccd1 vccd1 _19272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12716_ _12715_/X _12714_/X _12818_/S vssd1 vssd1 vccd1 vccd1 _12716_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13696_ _12638_/A _13665_/B _12639_/Y vssd1 vssd1 vccd1 vccd1 _13697_/B sky130_fd_sc_hd__o21ai_4
X_16484_ _10532_/B _19091_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _19091_/D sky130_fd_sc_hd__mux2_1
X_18223_ _19118_/CLK _18223_/D vssd1 vssd1 vccd1 vccd1 _18223_/Q sky130_fd_sc_hd__dfxtp_1
X_12647_ _13727_/A _12647_/B _13812_/A vssd1 vssd1 vccd1 vccd1 _12647_/Y sky130_fd_sc_hd__nor3_1
X_15435_ _18577_/Q _15465_/C _15434_/Y vssd1 vssd1 vccd1 vccd1 _15435_/X sky130_fd_sc_hd__a21o_1
XFILLER_248_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18154_ _19607_/CLK _18154_/D vssd1 vssd1 vccd1 vccd1 _18154_/Q sky130_fd_sc_hd__dfxtp_1
X_15366_ _15268_/B _15365_/X _15364_/Y vssd1 vssd1 vccd1 vccd1 _15368_/B sky130_fd_sc_hd__a21oi_1
X_12578_ _12578_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _12578_/Y sky130_fd_sc_hd__nor2_4
XFILLER_157_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ _19386_/Q _17115_/B vssd1 vssd1 vccd1 vccd1 _17105_/X sky130_fd_sc_hd__or2_1
X_14317_ _18174_/Q _17701_/A0 _14338_/S vssd1 vssd1 vccd1 vccd1 _18174_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11529_ _12626_/A _11678_/B _11293_/A vssd1 vssd1 vccd1 vccd1 _11677_/B sky130_fd_sc_hd__a21oi_4
X_18085_ _19304_/CLK _18085_/D vssd1 vssd1 vccd1 vccd1 _18085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15297_ _19465_/Q _19399_/Q vssd1 vssd1 vccd1 vccd1 _15299_/A sky130_fd_sc_hd__xnor2_1
XFILLER_171_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14248_ _18122_/Q _14266_/B vssd1 vssd1 vccd1 vccd1 _14248_/X sky130_fd_sc_hd__or2_1
X_17036_ _17199_/B _17046_/A2 _17035_/X _17106_/C1 vssd1 vssd1 vccd1 vccd1 _19354_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14179_ _14179_/A _14179_/B vssd1 vssd1 vccd1 vccd1 _18087_/D sky130_fd_sc_hd__and2_1
XFILLER_140_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout809 _14454_/Y vssd1 vssd1 vccd1 vccd1 _14486_/S sky130_fd_sc_hd__buf_12
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18987_ _19197_/CLK _18987_/D vssd1 vssd1 vccd1 vccd1 _18987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17938_ _18749_/CLK _17938_/D vssd1 vssd1 vccd1 vccd1 _17938_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1380 _11073_/B1 vssd1 vssd1 vccd1 vccd1 _11070_/S sky130_fd_sc_hd__buf_4
XFILLER_227_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1391 _10313_/S vssd1 vssd1 vccd1 vccd1 _10687_/S sky130_fd_sc_hd__buf_6
XFILLER_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17869_ _19310_/CLK _17869_/D vssd1 vssd1 vccd1 vccd1 _17869_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19608_ _19608_/CLK _19608_/D vssd1 vssd1 vccd1 vccd1 _19608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19539_ _19543_/CLK _19539_/D vssd1 vssd1 vccd1 vccd1 _19539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ _11046_/S1 _09217_/X _09220_/X _11053_/A vssd1 vssd1 vccd1 vccd1 _09223_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09154_ _09652_/A _09154_/B vssd1 vssd1 vccd1 vccd1 _09154_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _11706_/C _10027_/B vssd1 vssd1 vccd1 vccd1 _09085_/X sky130_fd_sc_hd__or2_1
XFILLER_206_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput90 dout0[52] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ _09987_/A _09987_/B vssd1 vssd1 vccd1 vccd1 _09987_/Y sky130_fd_sc_hd__nor2_1
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08938_ _08941_/B vssd1 vssd1 vccd1 vccd1 _08939_/C sky130_fd_sc_hd__inv_2
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ _17893_/Q _17892_/Q _09062_/B vssd1 vssd1 vccd1 vccd1 _12438_/B sky130_fd_sc_hd__nand3_2
XFILLER_123_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10900_ _10876_/Y _10880_/Y _11621_/C1 vssd1 vssd1 vccd1 vccd1 _10900_/X sky130_fd_sc_hd__a21o_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11880_ _11808_/X _11875_/A _11901_/B _11841_/X vssd1 vssd1 vccd1 vccd1 _11880_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10831_ _10831_/A vssd1 vssd1 vccd1 vccd1 _11537_/A sky130_fd_sc_hd__clkinv_2
XFILLER_26_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ _19251_/Q _13625_/A2 _13625_/B1 _19283_/Q vssd1 vssd1 vccd1 vccd1 _13550_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10762_ _19639_/Q _18928_/Q _11576_/S vssd1 vssd1 vccd1 vccd1 _10762_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12501_ _12501_/A _12501_/B vssd1 vssd1 vccd1 vccd1 _12553_/D sky130_fd_sc_hd__nand2_2
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13481_ _13541_/B _13481_/B vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__or2_1
XFILLER_9_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10693_ _18865_/Q _18897_/Q _11249_/S vssd1 vssd1 vccd1 vccd1 _10693_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15220_ _15263_/C vssd1 vssd1 vccd1 vccd1 _15220_/Y sky130_fd_sc_hd__inv_2
X_12432_ _11695_/B _12432_/A2 _09004_/X _12432_/B1 _18404_/Q vssd1 vssd1 vccd1 vccd1
+ _12433_/C sky130_fd_sc_hd__o32a_1
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15151_ _15151_/A _15259_/B vssd1 vssd1 vccd1 vccd1 _15151_/Y sky130_fd_sc_hd__nor2_1
X_12363_ _12429_/A1 _09652_/A _09329_/X _12417_/B1 _18381_/Q vssd1 vssd1 vccd1 vccd1
+ _12364_/B sky130_fd_sc_hd__o32ai_4
X_14102_ _17685_/A0 _18042_/Q _14106_/S vssd1 vssd1 vccd1 vccd1 _18042_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ _18453_/Q _18354_/Q _11325_/S vssd1 vssd1 vccd1 vccd1 _11314_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15082_ _15082_/A _15082_/B _15082_/C _12435_/A vssd1 vssd1 vccd1 vccd1 _15083_/B
+ sky130_fd_sc_hd__or4b_2
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12294_ _18085_/Q _12277_/B _14934_/C _18508_/Q vssd1 vssd1 vccd1 vccd1 _14672_/C
+ sky130_fd_sc_hd__a22o_2
XFILLER_153_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ _14033_/A1 _13886_/X _14032_/X _16153_/D vssd1 vssd1 vccd1 vccd1 _17981_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18910_ _19621_/CLK _18910_/D vssd1 vssd1 vccd1 vccd1 _18910_/Q sky130_fd_sc_hd__dfxtp_1
X_11245_ _11252_/S _11240_/X _11244_/X _11579_/A vssd1 vssd1 vccd1 vccd1 _11245_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_268_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18841_ _19628_/CLK _18841_/D vssd1 vssd1 vccd1 vccd1 _18841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _11155_/X _11158_/X _11175_/X vssd1 vssd1 vccd1 vccd1 _11176_/X sky130_fd_sc_hd__a21o_1
XFILLER_268_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10127_ _18046_/Q _18014_/Q _10206_/S vssd1 vssd1 vccd1 vccd1 _10127_/X sky130_fd_sc_hd__mux2_1
X_18772_ _18772_/CLK _18772_/D vssd1 vssd1 vccd1 vccd1 _18772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_283_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15984_ _18707_/Q _16016_/A2 _16147_/A2 _18756_/Q _16018_/C1 vssd1 vssd1 vccd1 vccd1
+ _15984_/X sky130_fd_sc_hd__a221o_1
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17723_ _17723_/A0 _19649_/Q _17723_/S vssd1 vssd1 vccd1 vccd1 _19649_/D sky130_fd_sc_hd__mux2_1
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10058_ _11274_/S1 _10047_/X _10057_/X _08950_/A vssd1 vssd1 vccd1 vccd1 _10058_/X
+ sky130_fd_sc_hd__o211a_1
X_14935_ _18125_/Q _14893_/S _14933_/X _14934_/X vssd1 vssd1 vccd1 vccd1 _14935_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17654_ _17720_/A0 _19582_/Q _17654_/S vssd1 vssd1 vccd1 vccd1 _19582_/D sky130_fd_sc_hd__mux2_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ input51/X input86/X _14947_/S vssd1 vssd1 vccd1 vccd1 _14867_/A sky130_fd_sc_hd__mux2_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16605_ _11376_/B _19208_/Q _16619_/S vssd1 vssd1 vccd1 vccd1 _19208_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13817_ _13810_/X _13813_/Y _13815_/Y _13816_/X vssd1 vssd1 vccd1 vccd1 _13817_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17585_ _17585_/A _17589_/B vssd1 vssd1 vccd1 vccd1 _17585_/X sky130_fd_sc_hd__or2_1
X_14797_ _14793_/Y _14796_/X _14950_/B1 vssd1 vssd1 vccd1 vccd1 _14797_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_69_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19630_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19324_ _19324_/CLK _19324_/D vssd1 vssd1 vccd1 vccd1 _19324_/Q sky130_fd_sc_hd__dfxtp_1
X_16536_ _17669_/A0 _19141_/Q _16556_/S vssd1 vssd1 vccd1 vccd1 _19141_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13748_ _19547_/Q _13946_/B vssd1 vssd1 vccd1 vccd1 _13748_/X sky130_fd_sc_hd__or2_1
XFILLER_250_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19255_ _19261_/CLK _19255_/D vssd1 vssd1 vccd1 vccd1 _19255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16467_ _16500_/A0 _19074_/Q _16488_/S vssd1 vssd1 vccd1 vccd1 _19074_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13679_ _13679_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13679_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18206_ _19133_/CLK _18206_/D vssd1 vssd1 vccd1 vccd1 _18206_/Q sky130_fd_sc_hd__dfxtp_1
X_15418_ _19470_/Q _19404_/Q vssd1 vssd1 vccd1 vccd1 _15419_/B sky130_fd_sc_hd__or2_1
XFILLER_192_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19186_ _19219_/CLK _19186_/D vssd1 vssd1 vccd1 vccd1 _19186_/Q sky130_fd_sc_hd__dfxtp_1
X_16398_ _16431_/A1 _19007_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _19007_/D sky130_fd_sc_hd__mux2_1
XFILLER_163_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18137_ _19138_/CLK _18137_/D vssd1 vssd1 vccd1 vccd1 _18137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15349_ _17129_/A _15348_/X _15424_/C1 vssd1 vssd1 vccd1 vccd1 _15349_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18068_ _19611_/CLK _18068_/D vssd1 vssd1 vccd1 vccd1 _18068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09910_ _09905_/X _09909_/Y _08947_/X vssd1 vssd1 vccd1 vccd1 _09910_/Y sky130_fd_sc_hd__a21oi_1
X_17019_ _19346_/Q _17041_/B vssd1 vssd1 vccd1 vccd1 _17019_/X sky130_fd_sc_hd__or2_1
XFILLER_171_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout606 _15080_/Y vssd1 vssd1 vccd1 vccd1 _17475_/A2 sky130_fd_sc_hd__buf_4
Xfanout617 _17557_/Y vssd1 vssd1 vccd1 vccd1 _17558_/B sky130_fd_sc_hd__buf_4
XFILLER_59_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09841_ _11252_/S _09834_/X _09840_/X vssd1 vssd1 vccd1 vccd1 _09859_/B sky130_fd_sc_hd__o21ai_2
Xfanout628 _16843_/X vssd1 vssd1 vccd1 vccd1 _16947_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_259_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout639 _17337_/S vssd1 vssd1 vccd1 vccd1 _17361_/S sky130_fd_sc_hd__buf_6
XFILLER_99_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09772_ _09752_/X _09754_/X _09771_/X _11252_/S _11579_/A vssd1 vssd1 vccd1 vccd1
+ _09772_/X sky130_fd_sc_hd__o221a_1
XFILLER_246_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09206_ _19628_/Q _18917_/Q _10128_/B vssd1 vssd1 vccd1 vccd1 _09206_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09137_ _09129_/X _09136_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09137_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _12756_/A _09080_/B _09068_/C _12261_/B vssd1 vssd1 vccd1 vccd1 _09083_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11030_ _11512_/A1 _18612_/Q _18183_/Q _11513_/B2 vssd1 vssd1 vccd1 vccd1 _11030_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12981_ _14214_/A _13028_/C vssd1 vssd1 vccd1 vccd1 _12982_/B sky130_fd_sc_hd__xnor2_4
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _14720_/A _14720_/B vssd1 vssd1 vccd1 vccd1 _14720_/Y sky130_fd_sc_hd__nor2_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11932_ _11939_/A1 _11822_/B _11935_/B1 input218/X vssd1 vssd1 vccd1 vccd1 _11932_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_273_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_500 _10364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_511 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_522 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14651_ _17710_/A0 _18457_/Q _14663_/S vssd1 vssd1 vccd1 vccd1 _18457_/D sky130_fd_sc_hd__mux2_1
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_533 _18396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _11899_/A _11863_/B _11863_/C vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__and3_4
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_544 _18109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _10810_/X _10811_/X _11606_/S vssd1 vssd1 vccd1 vccd1 _10814_/X sky130_fd_sc_hd__mux2_1
X_13602_ _13911_/A _13265_/Y _13266_/X _13602_/B2 vssd1 vssd1 vccd1 vccd1 _13602_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17370_ _17374_/A _17370_/B vssd1 vssd1 vccd1 vccd1 _19482_/D sky130_fd_sc_hd__and2_1
XFILLER_26_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11794_ _11820_/A _11820_/B vssd1 vssd1 vccd1 vccd1 _11794_/Y sky130_fd_sc_hd__nand2_1
X_14582_ _14592_/A _14582_/B vssd1 vssd1 vccd1 vccd1 _18399_/D sky130_fd_sc_hd__or2_1
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16321_ _17719_/A0 _18934_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _18934_/D sky130_fd_sc_hd__mux2_1
X_13533_ _13533_/A _13533_/B vssd1 vssd1 vccd1 vccd1 _14147_/B sky130_fd_sc_hd__xnor2_1
X_10745_ _10743_/X _10744_/X _10745_/S vssd1 vssd1 vccd1 vccd1 _10745_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19040_ _19653_/A _19040_/D vssd1 vssd1 vccd1 vccd1 _19040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16252_ _16418_/A0 _18867_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _18867_/D sky130_fd_sc_hd__mux2_1
X_13464_ _13476_/B _13961_/A vssd1 vssd1 vccd1 vccd1 _13464_/Y sky130_fd_sc_hd__nand2_1
XFILLER_199_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10676_ _10677_/A _12729_/A vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__nor2_4
XFILLER_199_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ _12427_/A _12415_/B vssd1 vssd1 vccd1 vccd1 _12415_/Y sky130_fd_sc_hd__nand2_1
X_15203_ _15189_/A _15186_/Y _15188_/B vssd1 vssd1 vccd1 vccd1 _15204_/B sky130_fd_sc_hd__o21ai_2
X_16183_ _16580_/A0 _18800_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _18800_/D sky130_fd_sc_hd__mux2_1
X_13395_ _13385_/Y _13388_/Y _13394_/X _12442_/C vssd1 vssd1 vccd1 vccd1 _13395_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12346_ _12349_/A _12346_/B vssd1 vssd1 vccd1 vccd1 _12346_/Y sky130_fd_sc_hd__nand2_1
X_15134_ _15216_/A1 _15131_/X _15786_/A2 _18103_/Q vssd1 vssd1 vccd1 vccd1 _15135_/B
+ sky130_fd_sc_hd__o2bb2a_2
Xclkbuf_leaf_187_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19611_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_116_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19291_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15065_ _18549_/Q _17676_/A0 _15079_/S vssd1 vssd1 vccd1 vccd1 _18549_/D sky130_fd_sc_hd__mux2_1
X_12277_ _12277_/A _12277_/B vssd1 vssd1 vccd1 vccd1 _12277_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14016_ _14036_/A _14016_/B vssd1 vssd1 vccd1 vccd1 _14016_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11228_ _11250_/A1 _18219_/Q _11154_/S _18954_/Q _11569_/S1 vssd1 vssd1 vccd1 vccd1
+ _11228_/X sky130_fd_sc_hd__o221a_1
XFILLER_141_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18824_ _19075_/CLK _18824_/D vssd1 vssd1 vccd1 vccd1 _18824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11159_ _18455_/Q _18356_/Q _11171_/S vssd1 vssd1 vccd1 vccd1 _11159_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18755_ _18761_/CLK _18755_/D vssd1 vssd1 vccd1 vccd1 _18755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15967_ _18699_/Q _15977_/A2 _15966_/X _14177_/A vssd1 vssd1 vccd1 vccd1 _18699_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput280 versionID[0] vssd1 vssd1 vccd1 vccd1 input280/X sky130_fd_sc_hd__buf_2
XFILLER_271_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17706_ _17706_/A0 _19632_/Q _17718_/S vssd1 vssd1 vccd1 vccd1 _19632_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14918_ _14979_/A1 _18271_/Q _14917_/Y _14918_/B1 vssd1 vssd1 vccd1 vccd1 _14918_/X
+ sky130_fd_sc_hd__a31o_1
X_18686_ _19276_/CLK _18686_/D vssd1 vssd1 vccd1 vccd1 _18686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15898_ _18675_/Q _15910_/A2 _15897_/X _15910_/C1 vssd1 vssd1 vccd1 vccd1 _18675_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17637_ _17703_/A0 _19565_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _19565_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14849_ _17806_/Q _15002_/B vssd1 vssd1 vccd1 vccd1 _14849_/X sky130_fd_sc_hd__or2_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17568_ _19526_/Q _17561_/B _17588_/B1 _17567_/X vssd1 vssd1 vccd1 vccd1 _19526_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19307_ _19326_/CLK _19307_/D vssd1 vssd1 vccd1 vccd1 _19307_/Q sky130_fd_sc_hd__dfxtp_1
X_16519_ _17685_/A0 _19125_/Q _16521_/S vssd1 vssd1 vccd1 vccd1 _19125_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17499_ _19511_/Q _17499_/A2 _17497_/X _17498_/Y _17360_/A vssd1 vssd1 vccd1 vccd1
+ _19511_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19238_ _19273_/CLK _19238_/D vssd1 vssd1 vccd1 vccd1 _19238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19169_ _19201_/CLK _19169_/D vssd1 vssd1 vccd1 vccd1 _19169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09824_ _11556_/C _09823_/X _09821_/X _11687_/A vssd1 vssd1 vccd1 vccd1 _09824_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_14__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_99_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09755_ _18535_/Q _18410_/Q _18019_/Q _17987_/Q _11073_/B1 _11559_/S1 vssd1 vssd1
+ vccd1 vccd1 _09755_/X sky130_fd_sc_hd__mux4_1
XFILLER_262_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_273_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09686_ _09683_/X _09685_/X _11484_/B1 vssd1 vssd1 vccd1 vccd1 _09686_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10530_ _10528_/X _10529_/X _08946_/B vssd1 vssd1 vccd1 vccd1 _10530_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10461_ _18464_/Q _18365_/Q _10613_/S vssd1 vssd1 vccd1 vccd1 _10461_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12200_ _17863_/Q _17864_/Q _12200_/C vssd1 vssd1 vccd1 vccd1 _12202_/B sky130_fd_sc_hd__and3_1
X_13180_ _13990_/B vssd1 vssd1 vccd1 vccd1 _13180_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10392_ _18262_/Q _18837_/Q _10864_/S vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12131_ _12219_/A _12136_/C vssd1 vssd1 vccd1 vccd1 _12131_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12062_ _17906_/Q _12086_/A2 _12061_/X _14340_/A vssd1 vssd1 vccd1 vccd1 _17808_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1902 _14991_/C1 vssd1 vssd1 vccd1 vccd1 _16787_/A sky130_fd_sc_hd__buf_6
XFILLER_150_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11013_ _18254_/Q _11395_/C _09129_/S _11012_/X vssd1 vssd1 vccd1 vccd1 _11013_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16870_ _17571_/A vssd1 vssd1 vccd1 vccd1 _16870_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout970 _14041_/Y vssd1 vssd1 vccd1 vccd1 _14064_/S sky130_fd_sc_hd__buf_6
Xfanout981 _12463_/X vssd1 vssd1 vccd1 vccd1 _13427_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _18613_/Q _17678_/A0 _15833_/S vssd1 vssd1 vccd1 vccd1 _18613_/D sky130_fd_sc_hd__mux2_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout992 _10531_/X vssd1 vssd1 vccd1 vccd1 _17716_/A0 sky130_fd_sc_hd__buf_4
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18540_ _19075_/CLK _18540_/D vssd1 vssd1 vccd1 vccd1 _18540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _19453_/Q _15793_/A2 _17208_/A vssd1 vssd1 vccd1 vccd1 _15752_/X sky130_fd_sc_hd__o21a_1
X_12964_ _15902_/A _12536_/Y _12505_/Y vssd1 vssd1 vccd1 vccd1 _12964_/X sky130_fd_sc_hd__a21o_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14703_ _17791_/Q _14702_/X _14993_/S vssd1 vssd1 vccd1 vccd1 _14703_/X sky130_fd_sc_hd__mux2_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18471_ _19229_/CLK _18471_/D vssd1 vssd1 vccd1 vccd1 _18471_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _18569_/Q _11918_/A2 _11706_/B _13125_/A vssd1 vssd1 vccd1 vccd1 _11915_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15683_ _15744_/A _15725_/A vssd1 vssd1 vccd1 vccd1 _15684_/B sky130_fd_sc_hd__and2_1
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12895_/A vssd1 vssd1 vccd1 vccd1 _12895_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_330 _11899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_341 _11482_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_352 _09086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17422_ _18107_/Q _17437_/A2 _17420_/X _17421_/X vssd1 vssd1 vccd1 vccd1 _17422_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_261_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14634_ _16593_/A0 _18440_/Q _14663_/S vssd1 vssd1 vccd1 vccd1 _18440_/D sky130_fd_sc_hd__mux2_1
XANTENNA_363 _12320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11846_ _11846_/A _11846_/B vssd1 vssd1 vccd1 vccd1 _11846_/Y sky130_fd_sc_hd__nand2_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_374 _18274_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_385 _17178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_396 _12599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _19474_/Q _17175_/B _17361_/S vssd1 vssd1 vccd1 vccd1 _17354_/B sky130_fd_sc_hd__mux2_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _11647_/A _11887_/B1 _11727_/B _11776_/Y vssd1 vssd1 vccd1 vccd1 _11777_/Y
+ sky130_fd_sc_hd__a211oi_4
X_14565_ _18391_/Q _14575_/A2 _14575_/B1 input19/X vssd1 vssd1 vccd1 vccd1 _14566_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16304_ _17702_/A0 _18917_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _18917_/D sky130_fd_sc_hd__mux2_1
X_13516_ _17841_/Q _13744_/A2 _13744_/B1 _17873_/Q vssd1 vssd1 vccd1 vccd1 _13516_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10728_ _10719_/S _10726_/X _10727_/X _11285_/S vssd1 vssd1 vccd1 vccd1 _10728_/X
+ sky130_fd_sc_hd__a211o_1
X_17284_ _19445_/Q _17313_/B _17283_/X vssd1 vssd1 vccd1 vccd1 _17285_/B sky130_fd_sc_hd__a21oi_1
XFILLER_201_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14496_ _17665_/A0 _18346_/Q _14517_/S vssd1 vssd1 vccd1 vccd1 _18346_/D sky130_fd_sc_hd__mux2_1
XFILLER_277_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19023_ _19055_/CLK _19023_/D vssd1 vssd1 vccd1 vccd1 _19023_/Q sky130_fd_sc_hd__dfxtp_1
X_16235_ _17699_/A0 _18850_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _18850_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ _17839_/Q _13744_/A2 _13744_/B1 _17871_/Q vssd1 vssd1 vccd1 vccd1 _13447_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10659_ _18617_/Q _18188_/Q _10667_/S vssd1 vssd1 vccd1 vccd1 _10659_/X sky130_fd_sc_hd__mux2_1
XFILLER_256_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13378_ _19310_/Q _12583_/Y _13376_/X _13377_/X vssd1 vssd1 vccd1 vccd1 _13378_/X
+ sky130_fd_sc_hd__a211o_1
X_16166_ _16431_/A1 _18783_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _18783_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15117_ _15117_/A _15123_/B vssd1 vssd1 vccd1 vccd1 _15118_/B sky130_fd_sc_hd__nor2_2
XFILLER_170_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12329_ _17821_/Q _17820_/Q _17819_/Q _17818_/Q vssd1 vssd1 vccd1 vccd1 _12330_/D
+ sky130_fd_sc_hd__or4bb_1
XFILLER_126_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16097_ _18751_/Q _16141_/B vssd1 vssd1 vccd1 vccd1 _16097_/Y sky130_fd_sc_hd__nand2_1
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15048_ _18532_/Q _16526_/A0 _15070_/S vssd1 vssd1 vccd1 vccd1 _18532_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18807_ _19646_/CLK _18807_/D vssd1 vssd1 vccd1 vccd1 _18807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16999_ _19336_/Q _17009_/B vssd1 vssd1 vccd1 vccd1 _16999_/X sky130_fd_sc_hd__or2_1
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09540_ _12471_/A0 _09539_/X _09538_/X vssd1 vssd1 vccd1 vccd1 _09540_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_84_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18817_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18738_ _18738_/CLK _18738_/D vssd1 vssd1 vccd1 vccd1 _18738_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19601_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09471_ _09469_/X _09470_/X _11024_/A1 vssd1 vssd1 vccd1 vccd1 _11800_/D sky130_fd_sc_hd__a21o_4
XFILLER_64_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18669_ _18715_/CLK _18669_/D vssd1 vssd1 vccd1 vccd1 _18669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1209 _12667_/X vssd1 vssd1 vccd1 vccd1 _12733_/S sky130_fd_sc_hd__buf_6
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09807_ _11284_/A1 _18207_/Q _11284_/B2 _18942_/Q _10040_/S vssd1 vssd1 vccd1 vccd1
+ _09807_/X sky130_fd_sc_hd__o221a_1
XFILLER_262_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09738_ input140/X input135/X _09990_/S vssd1 vssd1 vccd1 vccd1 _09738_/X sky130_fd_sc_hd__mux2_8
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09669_ _10689_/S _09669_/B vssd1 vssd1 vccd1 vccd1 _09669_/Y sky130_fd_sc_hd__nor2_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11700_ _18585_/Q _18584_/Q _18583_/Q _18582_/Q vssd1 vssd1 vccd1 vccd1 _11701_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_270_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12680_/A vssd1 vssd1 vccd1 vccd1 _12680_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _12656_/B _11631_/B vssd1 vssd1 vccd1 vccd1 _13958_/A sky130_fd_sc_hd__xnor2_4
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14350_ _14350_/A _16392_/C _14488_/C vssd1 vssd1 vccd1 vccd1 _16459_/C sky130_fd_sc_hd__or3_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11562_ _11560_/X _11561_/X _11562_/S vssd1 vssd1 vccd1 vccd1 _11562_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13301_ _19468_/Q _12529_/Y _12578_/Y _19340_/Q _13300_/X vssd1 vssd1 vccd1 vccd1
+ _13301_/X sky130_fd_sc_hd__a221o_1
X_10513_ _10511_/X _10512_/X _10513_/S vssd1 vssd1 vccd1 vccd1 _10513_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14281_ _17699_/A0 _18140_/Q _14304_/S vssd1 vssd1 vccd1 vccd1 _18140_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11493_ _11513_/A1 _18319_/Q _17770_/Q _10424_/S vssd1 vssd1 vccd1 vccd1 _11493_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16020_ _16020_/A _16056_/B vssd1 vssd1 vccd1 vccd1 _16020_/Y sky130_fd_sc_hd__nand2_2
X_13232_ _13136_/S _13042_/X _13197_/B1 vssd1 vssd1 vccd1 vccd1 _13232_/Y sky130_fd_sc_hd__o21bai_1
X_10444_ _11601_/A _10444_/B vssd1 vssd1 vccd1 vccd1 _10444_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13163_ _15259_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13163_/Y sky130_fd_sc_hd__nand2_1
X_10375_ _10368_/X _10374_/X _10358_/X vssd1 vssd1 vccd1 vccd1 _10375_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_152_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12114_ _17832_/Q _12114_/B vssd1 vssd1 vccd1 vccd1 _12120_/C sky130_fd_sc_hd__and2_2
XFILLER_124_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17971_ _18700_/CLK _17971_/D vssd1 vssd1 vccd1 vccd1 _17971_/Q sky130_fd_sc_hd__dfxtp_1
X_13094_ _13194_/S _13093_/Y _13197_/B1 vssd1 vssd1 vccd1 vccd1 _13094_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1710 _12488_/B vssd1 vssd1 vccd1 vccd1 _11406_/B2 sky130_fd_sc_hd__buf_12
X_16922_ _12482_/S _17939_/Q _16921_/X vssd1 vssd1 vccd1 vccd1 _17178_/B sky130_fd_sc_hd__o21a_4
X_12045_ _17800_/Q _12051_/B vssd1 vssd1 vccd1 vccd1 _12045_/X sky130_fd_sc_hd__or2_1
Xfanout1721 _18738_/Q vssd1 vssd1 vccd1 vccd1 _16034_/S sky130_fd_sc_hd__buf_6
XFILLER_266_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1732 _15088_/B vssd1 vssd1 vccd1 vccd1 _15092_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_278_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1743 _18273_/Q vssd1 vssd1 vccd1 vccd1 _14947_/S sky130_fd_sc_hd__buf_4
XFILLER_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19641_ _19641_/CLK _19641_/D vssd1 vssd1 vccd1 vccd1 _19641_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1754 _11252_/S vssd1 vssd1 vccd1 vccd1 _11583_/A sky130_fd_sc_hd__buf_12
Xfanout1765 _12466_/A0 vssd1 vssd1 vccd1 vccd1 _08843_/A sky130_fd_sc_hd__buf_12
X_16853_ _16852_/A _15837_/B _16852_/Y vssd1 vssd1 vccd1 vccd1 _17563_/A sky130_fd_sc_hd__o21ai_4
XFILLER_93_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1776 _17908_/Q vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__buf_12
XFILLER_281_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1787 _10513_/S vssd1 vssd1 vccd1 vccd1 _10663_/S sky130_fd_sc_hd__buf_8
XFILLER_253_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1798 _17822_/Q vssd1 vssd1 vccd1 vccd1 _08816_/A sky130_fd_sc_hd__buf_4
X_15804_ _18596_/Q _17661_/A0 _15817_/S vssd1 vssd1 vccd1 vccd1 _18596_/D sky130_fd_sc_hd__mux2_1
X_19572_ _19604_/CLK _19572_/D vssd1 vssd1 vccd1 vccd1 _19572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_265_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16784_ _16787_/A _16784_/B _16786_/B vssd1 vssd1 vccd1 vccd1 _19282_/D sky130_fd_sc_hd__nor3_1
XFILLER_219_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13996_ _14032_/B _13996_/B vssd1 vssd1 vccd1 vccd1 _13996_/Y sky130_fd_sc_hd__nand2_1
XFILLER_207_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18523_ _19286_/CLK _18523_/D vssd1 vssd1 vccd1 vccd1 _18523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15735_ _19484_/Q _19418_/Q vssd1 vssd1 vccd1 vccd1 _15756_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _13136_/S _12937_/Y _12946_/X vssd1 vssd1 vccd1 vccd1 _12947_/X sky130_fd_sc_hd__a21o_2
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18454_ _19640_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_1
X_15666_ _15789_/A1 _15665_/X _15789_/B1 vssd1 vssd1 vccd1 vccd1 _15666_/Y sky130_fd_sc_hd__a21oi_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _11972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ _12688_/X _12698_/X _12878_/S vssd1 vssd1 vccd1 vccd1 _12879_/B sky130_fd_sc_hd__mux2_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _13247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17405_ _19492_/Q _17423_/B _17403_/X _17404_/Y _17419_/C1 vssd1 vssd1 vccd1 vccd1
+ _19492_/D sky130_fd_sc_hd__o221a_1
XANTENNA_182 _14012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_193 _14028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14617_ _17676_/A0 _18424_/Q _14631_/S vssd1 vssd1 vccd1 vccd1 _18424_/D sky130_fd_sc_hd__mux2_1
X_11829_ _11865_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11829_/Y sky130_fd_sc_hd__nor2_2
X_18385_ _19471_/CLK _18385_/D vssd1 vssd1 vccd1 vccd1 _18385_/Q sky130_fd_sc_hd__dfxtp_4
X_15597_ _15787_/A _15639_/B vssd1 vssd1 vccd1 vccd1 _15620_/A sky130_fd_sc_hd__and2_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17336_ _17336_/A _17336_/B vssd1 vssd1 vccd1 vccd1 _19465_/D sky130_fd_sc_hd__and2_1
X_14548_ _14576_/A _14548_/B vssd1 vssd1 vccd1 vccd1 _18382_/D sky130_fd_sc_hd__or2_1
XFILLER_174_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_131_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19470_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17267_ _17265_/Y _17266_/X _17231_/A vssd1 vssd1 vccd1 vccd1 _19439_/D sky130_fd_sc_hd__a21oi_1
XFILLER_147_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14479_ _18331_/Q _17683_/A0 _14486_/S vssd1 vssd1 vccd1 vccd1 _18331_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19006_ _19589_/CLK _19006_/D vssd1 vssd1 vccd1 vccd1 _19006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16218_ _17715_/A0 _18834_/Q _16226_/S vssd1 vssd1 vccd1 vccd1 _18834_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17198_ _17198_/A _17198_/B vssd1 vssd1 vccd1 vccd1 _19417_/D sky130_fd_sc_hd__nor2_1
XFILLER_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16149_ _16149_/A _16149_/B vssd1 vssd1 vccd1 vccd1 _18774_/D sky130_fd_sc_hd__nor2_1
XFILLER_142_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08971_ _18637_/Q _18059_/Q _19078_/Q _18982_/Q _09306_/S _11510_/S1 vssd1 vssd1
+ vccd1 vccd1 _08972_/B sky130_fd_sc_hd__mux4_1
XFILLER_114_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09523_ _09523_/A _09523_/B _09523_/C vssd1 vssd1 vccd1 vccd1 _09523_/X sky130_fd_sc_hd__and3_2
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09454_ _09452_/X _09453_/X _09463_/S vssd1 vssd1 vccd1 vccd1 _09454_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09385_ _18540_/Q _18415_/Q _10128_/B vssd1 vssd1 vccd1 vccd1 _09385_/X sky130_fd_sc_hd__mux2_1
XFILLER_212_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10160_ _10160_/A _13913_/A vssd1 vssd1 vccd1 vccd1 _12656_/A sky130_fd_sc_hd__or2_4
XFILLER_105_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput370 _18372_/Q vssd1 vssd1 vccd1 vccd1 core_wb_stb_o sky130_fd_sc_hd__buf_4
Xoutput381 _11934_/X vssd1 vssd1 vccd1 vccd1 din0[14] sky130_fd_sc_hd__buf_4
Xfanout1006 _10081_/X vssd1 vssd1 vccd1 vccd1 _11489_/B1 sky130_fd_sc_hd__buf_4
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput392 _11944_/X vssd1 vssd1 vccd1 vccd1 din0[24] sky130_fd_sc_hd__buf_4
X_10091_ _19648_/Q _18937_/Q _10168_/S vssd1 vssd1 vccd1 vccd1 _10091_/X sky130_fd_sc_hd__mux2_1
Xfanout1017 _14402_/S vssd1 vssd1 vccd1 vccd1 _14412_/S sky130_fd_sc_hd__buf_12
XFILLER_273_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1028 _16530_/A0 vssd1 vssd1 vccd1 vccd1 _17663_/A0 sky130_fd_sc_hd__buf_2
XFILLER_102_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1039 _11488_/A vssd1 vssd1 vccd1 vccd1 _11103_/A sky130_fd_sc_hd__buf_4
XFILLER_248_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13850_ _19420_/Q _13948_/A2 _13948_/B1 vssd1 vssd1 vccd1 vccd1 _13850_/X sky130_fd_sc_hd__a21o_1
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12801_ _12676_/X _12681_/X _12823_/A vssd1 vssd1 vccd1 vccd1 _12938_/B sky130_fd_sc_hd__mux2_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10993_ _10403_/S _10992_/X _10991_/X _11478_/S vssd1 vssd1 vccd1 vccd1 _10993_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_262_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13781_ _19516_/Q _13781_/A2 _13781_/B1 _13780_/X vssd1 vssd1 vccd1 vccd1 _13781_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15520_ _19474_/Q _19408_/Q vssd1 vssd1 vccd1 vccd1 _15521_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12598_/A _12641_/B _12732_/S vssd1 vssd1 vccd1 vccd1 _12821_/B sky130_fd_sc_hd__mux2_2
XFILLER_203_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _15502_/B _13473_/Y _15133_/B _15450_/Y vssd1 vssd1 vccd1 vccd1 _15452_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _11627_/Y _12663_/B vssd1 vssd1 vccd1 vccd1 _14156_/S sky130_fd_sc_hd__nand2b_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14402_ _17709_/A0 _18253_/Q _14402_/S vssd1 vssd1 vccd1 vccd1 _18253_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18170_ _18880_/CLK _18170_/D vssd1 vssd1 vccd1 vccd1 _18170_/Q sky130_fd_sc_hd__dfxtp_1
X_11614_ _18657_/Q _18079_/Q _11617_/S vssd1 vssd1 vccd1 vccd1 _11614_/X sky130_fd_sc_hd__mux2_1
X_15382_ _18114_/Q _15133_/Y _15381_/X _15382_/B2 vssd1 vssd1 vccd1 vccd1 _15387_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12594_/A _12594_/B vssd1 vssd1 vccd1 vccd1 _12594_/X sky130_fd_sc_hd__or2_1
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ _15119_/Y _17394_/A _17120_/Y _17141_/A vssd1 vssd1 vccd1 vccd1 _17121_/X
+ sky130_fd_sc_hd__a31o_1
X_14333_ _18190_/Q _17717_/A0 _14339_/S vssd1 vssd1 vccd1 vccd1 _18190_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11545_ _11545_/A _11545_/B vssd1 vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__nor2_4
XFILLER_7_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17052_ _17052_/A _17052_/B _17052_/C _17052_/D vssd1 vssd1 vccd1 vccd1 _17316_/B
+ sky130_fd_sc_hd__or4_4
X_11476_ _18248_/Q _18823_/Q _11477_/S vssd1 vssd1 vccd1 vccd1 _11476_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14264_ _18130_/Q _14266_/B vssd1 vssd1 vccd1 vccd1 _14264_/X sky130_fd_sc_hd__or2_1
XFILLER_125_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16003_ _18717_/Q _16003_/A2 _16002_/X _14205_/A vssd1 vssd1 vccd1 vccd1 _18717_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10427_ _11506_/A1 _18230_/Q _10424_/S _18965_/Q _10427_/C1 vssd1 vssd1 vccd1 vccd1
+ _10427_/X sky130_fd_sc_hd__o221a_1
X_13215_ _17864_/Q _13945_/A2 _13207_/X _13945_/B2 _13952_/B1 vssd1 vssd1 vccd1 vccd1
+ _13215_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ _14197_/A _14195_/B vssd1 vssd1 vccd1 vccd1 _18095_/D sky130_fd_sc_hd__and2_1
XFILLER_83_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10358_ _11053_/A _10352_/X _10355_/X _10357_/X _11417_/B1 vssd1 vssd1 vccd1 vccd1
+ _10358_/X sky130_fd_sc_hd__a311o_4
XFILLER_97_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13146_ _13257_/A _13146_/B vssd1 vssd1 vccd1 vccd1 _17927_/D sky130_fd_sc_hd__and2_1
XFILLER_151_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17954_ _17958_/CLK _17954_/D vssd1 vssd1 vccd1 vccd1 _17954_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13077_ _13757_/A _13986_/B _13058_/X vssd1 vssd1 vccd1 vccd1 _13079_/B sky130_fd_sc_hd__o21ai_1
X_10289_ _18264_/Q _18839_/Q _10299_/S vssd1 vssd1 vccd1 vccd1 _10289_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16905_ _18757_/Q _16961_/A2 _16969_/B1 input221/X _16969_/C1 vssd1 vssd1 vccd1 vccd1
+ _16905_/X sky130_fd_sc_hd__a221o_2
Xfanout1540 _10653_/A1 vssd1 vssd1 vccd1 vccd1 _09967_/S sky130_fd_sc_hd__buf_8
X_12028_ _17889_/Q _12035_/B _12027_/X _12350_/C1 vssd1 vssd1 vccd1 vccd1 _17791_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1551 _10280_/S vssd1 vssd1 vccd1 vccd1 _10371_/S sky130_fd_sc_hd__buf_8
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17885_ _19327_/CLK _17885_/D vssd1 vssd1 vccd1 vccd1 _17885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1562 _08898_/Y vssd1 vssd1 vccd1 vccd1 _11286_/B1 sky130_fd_sc_hd__buf_12
XFILLER_238_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1573 fanout1581/X vssd1 vssd1 vccd1 vccd1 _10653_/C1 sky130_fd_sc_hd__buf_6
Xfanout1584 _10211_/A1 vssd1 vssd1 vccd1 vccd1 _10881_/S1 sky130_fd_sc_hd__buf_6
XFILLER_253_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1595 _08904_/A vssd1 vssd1 vccd1 vccd1 _11053_/A sky130_fd_sc_hd__clkbuf_16
X_19624_ _19624_/CLK _19624_/D vssd1 vssd1 vccd1 vccd1 _19624_/Q sky130_fd_sc_hd__dfxtp_1
X_16836_ _17821_/Q _12285_/A _16836_/S vssd1 vssd1 vccd1 vccd1 _17052_/B sky130_fd_sc_hd__mux2_1
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19555_ _19587_/CLK _19555_/D vssd1 vssd1 vccd1 vccd1 _19555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16767_ _19276_/Q _19275_/Q _16767_/C vssd1 vssd1 vccd1 vccd1 _16770_/B sky130_fd_sc_hd__and3_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13979_ _17954_/Q _14004_/A _13978_/Y _13981_/C1 vssd1 vssd1 vccd1 vccd1 _17954_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18506_ _19229_/CLK _18506_/D vssd1 vssd1 vccd1 vccd1 _18506_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_207_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15718_ _18589_/Q _15718_/A2 _15717_/X _15718_/C1 vssd1 vssd1 vccd1 vccd1 _18589_/D
+ sky130_fd_sc_hd__o211a_1
X_19486_ _19522_/CLK _19486_/D vssd1 vssd1 vccd1 vccd1 _19486_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16698_ _16795_/A _16704_/C vssd1 vssd1 vccd1 vccd1 _16698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18437_ _19225_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_278_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15649_ _19480_/Q _19414_/Q vssd1 vssd1 vccd1 vccd1 _15651_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09170_ _18026_/Q _17994_/Q _09181_/S vssd1 vssd1 vccd1 vccd1 _09170_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18368_ _19646_/CLK _18368_/D vssd1 vssd1 vccd1 vccd1 _18368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17319_ _19457_/Q _17123_/B _17345_/S vssd1 vssd1 vccd1 vccd1 _17320_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18299_ _19448_/CLK _18299_/D vssd1 vssd1 vccd1 vccd1 _18299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput109 dout1[11] vssd1 vssd1 vccd1 vccd1 input109/X sky130_fd_sc_hd__clkbuf_2
X_08954_ _08954_/A _08956_/C _08954_/C vssd1 vssd1 vccd1 vccd1 _09055_/C sky130_fd_sc_hd__and3_1
XFILLER_257_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08885_ _18593_/Q _18592_/Q _18591_/Q vssd1 vssd1 vccd1 vccd1 _11724_/B sky130_fd_sc_hd__or3_4
XFILLER_257_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09506_ _09504_/X _09505_/X _10373_/S vssd1 vssd1 vccd1 vccd1 _09506_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _09859_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _11800_/C sky130_fd_sc_hd__or2_2
XFILLER_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09368_ _19043_/Q _19011_/Q _10141_/S vssd1 vssd1 vccd1 vccd1 _09368_/X sky130_fd_sc_hd__mux2_1
X_09299_ _18541_/Q _18416_/Q _09306_/S vssd1 vssd1 vccd1 vccd1 _09299_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_60 _10121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _11310_/X _11313_/X _11329_/X vssd1 vssd1 vccd1 vccd1 _11330_/X sky130_fd_sc_hd__a21o_1
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_93 _10837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11261_ _18116_/Q _11337_/B vssd1 vssd1 vccd1 vccd1 _11261_/X sky130_fd_sc_hd__or2_2
XFILLER_273_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10212_ _19064_/Q _19032_/Q _10215_/S vssd1 vssd1 vccd1 vccd1 _10212_/X sky130_fd_sc_hd__mux2_1
X_13000_ _13912_/B1 _12999_/X _09736_/B vssd1 vssd1 vccd1 vccd1 _13000_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_268_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11192_ _11190_/X _11191_/X _11198_/S vssd1 vssd1 vccd1 vccd1 _11192_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10143_ _18905_/Q _10217_/B vssd1 vssd1 vccd1 vccd1 _10143_/X sky130_fd_sc_hd__or2_1
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ _18496_/Q _15011_/A2 _14950_/Y _16787_/A vssd1 vssd1 vccd1 vccd1 _18496_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10074_ _11742_/B _10074_/B vssd1 vssd1 vccd1 vccd1 _11746_/A sky130_fd_sc_hd__nand2_2
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13902_ _13934_/B _13902_/B vssd1 vssd1 vccd1 vccd1 _13903_/B sky130_fd_sc_hd__nor2_2
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17670_ _17670_/A0 _19597_/Q _17689_/S vssd1 vssd1 vccd1 vccd1 _19597_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14882_ _17809_/Q _15002_/B _14881_/X vssd1 vssd1 vccd1 vccd1 _14882_/X sky130_fd_sc_hd__o21a_1
XFILLER_247_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16621_ _16621_/A0 _19224_/Q _16622_/S vssd1 vssd1 vccd1 vccd1 _19224_/D sky130_fd_sc_hd__mux2_1
X_13833_ _13758_/A _13818_/X _13956_/B1 vssd1 vssd1 vccd1 vccd1 _13833_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19340_ _19502_/CLK _19340_/D vssd1 vssd1 vccd1 vccd1 _19340_/Q sky130_fd_sc_hd__dfxtp_1
X_16552_ _17685_/A0 _19157_/Q _16554_/S vssd1 vssd1 vccd1 vccd1 _19157_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13764_ _13761_/B _14150_/A _13892_/B1 vssd1 vssd1 vccd1 vccd1 _13764_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _10952_/Y _10956_/Y _11621_/C1 vssd1 vssd1 vccd1 vccd1 _10976_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15503_ _15526_/B _13542_/X _15133_/B _15502_/Y vssd1 vssd1 vccd1 vccd1 _15503_/X
+ sky130_fd_sc_hd__a31o_1
X_19271_ _19273_/CLK _19271_/D vssd1 vssd1 vccd1 vccd1 _19271_/Q sky130_fd_sc_hd__dfxtp_1
X_12715_ _12613_/B _12649_/B _12733_/S vssd1 vssd1 vccd1 vccd1 _12715_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16483_ _16549_/A0 _19090_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _19090_/D sky130_fd_sc_hd__mux2_1
XFILLER_241_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13695_ _13695_/A _13761_/B vssd1 vssd1 vccd1 vccd1 _13695_/X sky130_fd_sc_hd__or2_1
XFILLER_231_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18222_ _19604_/CLK _18222_/D vssd1 vssd1 vccd1 vccd1 _18222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15434_ _18577_/Q _15465_/C _15437_/B1 vssd1 vssd1 vccd1 vccd1 _15434_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_175_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12646_ _13597_/B _12638_/Y _12645_/X vssd1 vssd1 vccd1 vccd1 _13727_/B sky130_fd_sc_hd__a21o_4
XFILLER_62_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18153_ _19607_/CLK _18153_/D vssd1 vssd1 vccd1 vccd1 _18153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15365_ _15365_/A _15365_/B _15365_/C _15365_/D vssd1 vssd1 vccd1 vccd1 _15365_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_178_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12577_ _12577_/A _12577_/B vssd1 vssd1 vccd1 vccd1 _12582_/B sky130_fd_sc_hd__or2_4
XFILLER_156_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17104_ _17196_/B _17116_/A2 _17103_/X _17368_/A vssd1 vssd1 vccd1 vccd1 _19385_/D
+ sky130_fd_sc_hd__o211a_1
X_14316_ _18173_/Q _17700_/A0 _14335_/S vssd1 vssd1 vccd1 vccd1 _18173_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18084_ _19304_/CLK _18084_/D vssd1 vssd1 vccd1 vccd1 _18084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11528_ _13387_/A _11679_/B _11369_/A vssd1 vssd1 vccd1 vccd1 _11678_/B sky130_fd_sc_hd__o21bai_4
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15296_ _19433_/Q _15411_/B _17166_/A _15295_/X vssd1 vssd1 vccd1 vccd1 _15296_/X
+ sky130_fd_sc_hd__o211a_1
X_17035_ _19354_/Q _17041_/B vssd1 vssd1 vccd1 vccd1 _17035_/X sky130_fd_sc_hd__or2_1
X_14247_ _18295_/Q _14247_/A2 _14246_/X _14442_/B vssd1 vssd1 vccd1 vccd1 _18121_/D
+ sky130_fd_sc_hd__o211a_1
X_11459_ _11459_/A1 _11457_/X _11458_/X _11459_/B1 vssd1 vssd1 vccd1 vccd1 _11459_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_264_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14178_ _18700_/Q _18087_/Q _14186_/S vssd1 vssd1 vccd1 vccd1 _14179_/B sky130_fd_sc_hd__mux2_1
XFILLER_113_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13129_ _13130_/A _13129_/B vssd1 vssd1 vccd1 vccd1 _13129_/Y sky130_fd_sc_hd__nor2_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _19146_/CLK _18986_/D vssd1 vssd1 vccd1 vccd1 _18986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17937_ _18700_/CLK _17937_/D vssd1 vssd1 vccd1 vccd1 _17937_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1370 _10856_/C vssd1 vssd1 vccd1 vccd1 _10929_/S sky130_fd_sc_hd__buf_4
XFILLER_239_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17868_ _19327_/CLK _17868_/D vssd1 vssd1 vccd1 vccd1 _17868_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1381 fanout1386/X vssd1 vssd1 vccd1 vccd1 _11073_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout1392 _10320_/S vssd1 vssd1 vccd1 vccd1 _10313_/S sky130_fd_sc_hd__buf_6
XFILLER_26_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19607_ _19607_/CLK _19607_/D vssd1 vssd1 vccd1 vccd1 _19607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16819_ _16819_/A _16819_/B _16819_/C vssd1 vssd1 vccd1 vccd1 _16819_/Y sky130_fd_sc_hd__nor3_1
X_17799_ _17930_/CLK _17799_/D vssd1 vssd1 vccd1 vccd1 _17799_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_254_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19538_ _19543_/CLK _19538_/D vssd1 vssd1 vccd1 vccd1 _19538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19469_ _19502_/CLK _19469_/D vssd1 vssd1 vccd1 vccd1 _19469_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09222_ _11046_/S1 _09212_/X _09221_/X _11438_/B1 vssd1 vssd1 vccd1 vccd1 _09222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09153_ input108/X input143/X _09651_/S vssd1 vssd1 vccd1 vccd1 _09154_/B sky130_fd_sc_hd__mux2_4
XFILLER_159_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09084_ _11706_/C _10027_/B vssd1 vssd1 vccd1 vccd1 _09140_/S sky130_fd_sc_hd__nor2_4
XFILLER_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput80 dout0[43] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput91 dout0[53] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ _11217_/A _09986_/B _09986_/C vssd1 vssd1 vccd1 vccd1 _09987_/B sky130_fd_sc_hd__and3_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08937_ _08991_/A _17796_/Q _17794_/Q vssd1 vssd1 vccd1 vccd1 _08941_/B sky130_fd_sc_hd__or3b_2
XFILLER_218_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08868_ _17892_/Q _09062_/B vssd1 vssd1 vccd1 vccd1 _09070_/D sky130_fd_sc_hd__nand2_2
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10830_ _10832_/A _12640_/B vssd1 vssd1 vccd1 vccd1 _10831_/A sky130_fd_sc_hd__or2_2
XFILLER_60_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _18460_/Q _18361_/Q _11576_/S vssd1 vssd1 vccd1 vccd1 _10761_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12500_ _12577_/A _12582_/A vssd1 vssd1 vccd1 vccd1 _13167_/A sky130_fd_sc_hd__or2_4
XFILLER_279_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10692_ _10690_/X _10691_/X _11248_/S vssd1 vssd1 vccd1 vccd1 _10692_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13480_ _14238_/A _13479_/C _18118_/Q vssd1 vssd1 vccd1 vccd1 _13481_/B sky130_fd_sc_hd__a21oi_1
XFILLER_232_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12431_ _12442_/A _12430_/A _12430_/Y _14001_/C1 vssd1 vssd1 vccd1 vccd1 _17918_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15150_ _08852_/Y _15381_/A3 _12761_/B _09777_/A vssd1 vssd1 vccd1 vccd1 _15155_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_12362_ _17887_/Q _12433_/B _12361_/X _12360_/X _12383_/C1 vssd1 vssd1 vccd1 vccd1
+ _17895_/D sky130_fd_sc_hd__o311a_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14101_ _16551_/A0 _18041_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _18041_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11313_ _10785_/A _11311_/X _11312_/X _11563_/B1 vssd1 vssd1 vccd1 vccd1 _11313_/X
+ sky130_fd_sc_hd__o31a_1
X_12293_ _18086_/Q _12277_/B _14934_/C _18509_/Q vssd1 vssd1 vccd1 vccd1 _14680_/B
+ sky130_fd_sc_hd__a22o_2
X_15081_ _15081_/A _15120_/B vssd1 vssd1 vccd1 vccd1 _17531_/B sky130_fd_sc_hd__or2_2
X_14032_ _17981_/Q _14032_/B vssd1 vssd1 vccd1 vccd1 _14032_/X sky130_fd_sc_hd__or2_1
X_11244_ _09095_/A _11241_/X _11242_/X _11243_/X vssd1 vssd1 vccd1 vccd1 _11244_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18840_ _19225_/CLK _18840_/D vssd1 vssd1 vccd1 vccd1 _18840_/Q sky130_fd_sc_hd__dfxtp_1
X_11175_ _11148_/X _11151_/X _10326_/A vssd1 vssd1 vccd1 vccd1 _11175_/X sky130_fd_sc_hd__a21o_1
XFILLER_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10126_ _10219_/A1 _19584_/Q _10206_/S _19616_/Q _10205_/S vssd1 vssd1 vccd1 vccd1
+ _10126_/X sky130_fd_sc_hd__o221a_1
X_18771_ _18775_/CLK _18771_/D vssd1 vssd1 vccd1 vccd1 _18771_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15983_ _18707_/Q _16005_/A2 _15982_/X _16972_/A vssd1 vssd1 vccd1 vccd1 _18707_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ _17722_/A0 _19648_/Q _17722_/S vssd1 vssd1 vccd1 vccd1 _19648_/D sky130_fd_sc_hd__mux2_1
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14934_ _19230_/Q _15014_/B _14934_/C _14934_/D vssd1 vssd1 vccd1 vccd1 _14934_/X
+ sky130_fd_sc_hd__and4_4
X_10057_ _10719_/S _10049_/X _10048_/X _11198_/S vssd1 vssd1 vccd1 vccd1 _10057_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17653_ _17686_/A0 _19581_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _19581_/D sky130_fd_sc_hd__mux2_1
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ _14865_/A1 _14864_/X _14865_/B1 vssd1 vssd1 vccd1 vccd1 _14865_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16604_ _11452_/B _19207_/Q _16619_/S vssd1 vssd1 vccd1 vccd1 _19207_/D sky130_fd_sc_hd__mux2_1
XFILLER_263_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13816_ _12704_/S _12998_/X _13002_/X _13863_/B2 vssd1 vssd1 vccd1 vccd1 _13816_/X
+ sky130_fd_sc_hd__o22a_1
X_17584_ _19534_/Q _17558_/B _17603_/B1 _17583_/X vssd1 vssd1 vccd1 vccd1 _19534_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_250_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14796_ _14696_/A _18270_/Q _14795_/Y _14846_/B1 vssd1 vssd1 vccd1 vccd1 _14796_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_63_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19323_ _19323_/CLK _19323_/D vssd1 vssd1 vccd1 vccd1 _19323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16535_ _16535_/A0 _19140_/Q _16556_/S vssd1 vssd1 vccd1 vccd1 _19140_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13747_ _17880_/Q _13747_/A2 _13745_/X _13747_/B2 _13854_/B1 vssd1 vssd1 vccd1 vccd1
+ _13747_/X sky130_fd_sc_hd__a221o_1
X_10959_ _11594_/A1 _18958_/Q _18223_/Q _11125_/B2 vssd1 vssd1 vccd1 vccd1 _10959_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19254_ _19261_/CLK _19254_/D vssd1 vssd1 vccd1 vccd1 _19254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16466_ _16532_/A0 _19073_/Q _16485_/S vssd1 vssd1 vccd1 vccd1 _19073_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13678_ _17942_/Q _13973_/A2 _13677_/X _14417_/A vssd1 vssd1 vccd1 vccd1 _17942_/D
+ sky130_fd_sc_hd__o211a_1
X_18205_ _19201_/CLK _18205_/D vssd1 vssd1 vccd1 vccd1 _18205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15417_ _19470_/Q _19404_/Q vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__nand2_1
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19185_ _19623_/CLK _19185_/D vssd1 vssd1 vccd1 vccd1 _19185_/Q sky130_fd_sc_hd__dfxtp_1
X_12629_ _12597_/Y _12628_/X _13411_/A _13387_/A vssd1 vssd1 vccd1 vccd1 _12629_/X
+ sky130_fd_sc_hd__o211a_1
X_16397_ _16595_/A0 _19006_/Q _16425_/S vssd1 vssd1 vccd1 vccd1 _19006_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19591_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18136_ _19589_/CLK _18136_/D vssd1 vssd1 vccd1 vccd1 _18136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15348_ _19467_/Q _15347_/Y _15498_/S vssd1 vssd1 vccd1 vccd1 _15348_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18067_ _19118_/CLK _18067_/D vssd1 vssd1 vccd1 vccd1 _18067_/Q sky130_fd_sc_hd__dfxtp_1
X_15279_ _19463_/Q _19397_/Q _15278_/X vssd1 vssd1 vccd1 vccd1 _15280_/B sky130_fd_sc_hd__o21ai_4
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17018_ _17172_/B _17032_/A2 _17017_/X _17352_/A vssd1 vssd1 vccd1 vccd1 _19345_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout607 _13951_/C1 vssd1 vssd1 vccd1 vccd1 _13884_/C1 sky130_fd_sc_hd__buf_8
X_09840_ _09750_/S _09839_/X _10326_/A vssd1 vssd1 vccd1 vccd1 _09840_/X sky130_fd_sc_hd__o21a_1
Xfanout618 _17120_/B vssd1 vssd1 vccd1 vccd1 _17119_/B sky130_fd_sc_hd__buf_4
Xfanout629 _16843_/X vssd1 vssd1 vccd1 vccd1 _16971_/S sky130_fd_sc_hd__buf_6
XFILLER_59_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_13__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_09771_ _09769_/X _09770_/X _11084_/S vssd1 vssd1 vccd1 vccd1 _09771_/X sky130_fd_sc_hd__mux2_1
X_18969_ _19225_/CLK _18969_/D vssd1 vssd1 vccd1 vccd1 _18969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09205_ _18449_/Q _18350_/Q _10128_/B vssd1 vssd1 vccd1 vccd1 _09205_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09136_ _09133_/X _09135_/X _09136_/S vssd1 vssd1 vccd1 vccd1 _09136_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ _17894_/Q _12443_/A vssd1 vssd1 vccd1 vccd1 _09068_/C sky130_fd_sc_hd__or2_1
XFILLER_118_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09969_ _18017_/Q _17985_/Q _09973_/S vssd1 vssd1 vccd1 vccd1 _09969_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12980_ _13930_/A1 _12962_/X _13253_/B1 vssd1 vssd1 vccd1 vccd1 _12980_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_217_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11931_ _11810_/A _11944_/A1 _11818_/C _11959_/A2 input217/X vssd1 vssd1 vccd1 vccd1
+ _11931_/X sky130_fd_sc_hd__a32o_4
XFILLER_100_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_501 _12320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_512 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_523 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14650_ _17709_/A0 _18456_/Q _14664_/S vssd1 vssd1 vccd1 vccd1 _18456_/D sky130_fd_sc_hd__mux2_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11862_ _11846_/A _11826_/A _11825_/B _11861_/Y vssd1 vssd1 vccd1 vccd1 _11863_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_534 _15854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_545 _12073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13601_ _13962_/B _13600_/X _10909_/B vssd1 vssd1 vccd1 vccd1 _13601_/X sky130_fd_sc_hd__a21o_1
XFILLER_261_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10813_ _11360_/A1 _19216_/Q _19184_/Q _11360_/B2 _08899_/A vssd1 vssd1 vccd1 vccd1
+ _10813_/X sky130_fd_sc_hd__a221o_1
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _18399_/Q _14589_/A2 _14589_/B1 input28/X vssd1 vssd1 vccd1 vccd1 _14582_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_260_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11793_ _11816_/A _11793_/B vssd1 vssd1 vccd1 vccd1 _11820_/B sky130_fd_sc_hd__nor2_8
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16320_ _17718_/A0 _18933_/Q _16320_/S vssd1 vssd1 vccd1 vccd1 _18933_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13532_ _11676_/A _13466_/A _12632_/X vssd1 vssd1 vccd1 vccd1 _13533_/B sky130_fd_sc_hd__a21boi_2
XFILLER_185_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10744_ _19640_/Q _18929_/Q _10744_/S vssd1 vssd1 vccd1 vccd1 _10744_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16251_ _17715_/A0 _18866_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _18866_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ _13622_/A _13476_/B _13323_/X _13462_/X vssd1 vssd1 vccd1 vccd1 _13463_/X
+ sky130_fd_sc_hd__a211o_1
X_10675_ _12729_/A vssd1 vssd1 vccd1 vccd1 _10675_/Y sky130_fd_sc_hd__inv_2
X_15202_ _19461_/Q _19395_/Q vssd1 vssd1 vccd1 vccd1 _15204_/A sky130_fd_sc_hd__xnor2_1
X_12414_ _18398_/Q _12429_/B1 _09232_/Y _08858_/A vssd1 vssd1 vccd1 vccd1 _12415_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_185_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16182_ _17712_/A0 _18799_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _18799_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13394_ _13863_/B2 _13390_/X _13391_/Y _12704_/S _13393_/X vssd1 vssd1 vccd1 vccd1
+ _13394_/X sky130_fd_sc_hd__o221a_1
XFILLER_126_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15133_ _15133_/A _15133_/B vssd1 vssd1 vccd1 vccd1 _15133_/Y sky130_fd_sc_hd__nand2_8
X_12345_ _11695_/B _09991_/A _09822_/X _12432_/B1 _18375_/Q vssd1 vssd1 vccd1 vccd1
+ _12346_/B sky130_fd_sc_hd__o32ai_4
XFILLER_141_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15064_ _18548_/Q _17708_/A0 _15070_/S vssd1 vssd1 vccd1 vccd1 _18548_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12276_ _12276_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _12276_/X sky130_fd_sc_hd__or2_2
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14015_ _17972_/Q _14036_/A _14014_/Y _14037_/C1 vssd1 vssd1 vccd1 vccd1 _17972_/D
+ sky130_fd_sc_hd__o211a_1
X_11227_ _11567_/S _11226_/X _11225_/X _11248_/S vssd1 vssd1 vccd1 vccd1 _11227_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_268_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18823_ _18884_/CLK _18823_/D vssd1 vssd1 vccd1 vccd1 _18823_/Q sky130_fd_sc_hd__dfxtp_1
X_11158_ _10707_/A _11156_/X _11157_/X _11237_/B1 vssd1 vssd1 vccd1 vccd1 _11158_/X
+ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_156_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19471_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_283_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10109_ _10107_/X _10108_/X _10335_/S vssd1 vssd1 vccd1 vccd1 _10109_/X sky130_fd_sc_hd__mux2_1
X_18754_ _18776_/CLK _18754_/D vssd1 vssd1 vccd1 vccd1 _18754_/Q sky130_fd_sc_hd__dfxtp_1
X_15966_ _18698_/Q _15970_/A2 _15976_/B1 _18747_/Q _15976_/C1 vssd1 vssd1 vccd1 vccd1
+ _15966_/X sky130_fd_sc_hd__a221o_1
X_11089_ _11583_/A _11084_/X _11088_/X _11579_/A vssd1 vssd1 vccd1 vccd1 _11089_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput270 partID[15] vssd1 vssd1 vccd1 vccd1 input270/X sky130_fd_sc_hd__clkbuf_4
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput281 versionID[1] vssd1 vssd1 vccd1 vccd1 _12770_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17705_ _17705_/A0 _19631_/Q _17722_/S vssd1 vssd1 vccd1 vccd1 _19631_/D sky130_fd_sc_hd__mux2_1
X_14917_ _14917_/A vssd1 vssd1 vccd1 vccd1 _14917_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_64_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18685_ _19276_/CLK _18685_/D vssd1 vssd1 vccd1 vccd1 _18685_/Q sky130_fd_sc_hd__dfxtp_1
X_15897_ _18674_/Q _15906_/A2 _15905_/C _15896_/Y _15903_/B1 vssd1 vssd1 vccd1 vccd1
+ _15897_/X sky130_fd_sc_hd__a221o_1
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17636_ _17669_/A0 _19564_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _19564_/D sky130_fd_sc_hd__mux2_1
XFILLER_223_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14848_ _18486_/Q _15001_/A2 _14847_/Y _16808_/A vssd1 vssd1 vccd1 vccd1 _18486_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17567_ _17567_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17567_/X sky130_fd_sc_hd__or2_1
X_14779_ _16392_/B _14982_/B vssd1 vssd1 vccd1 vccd1 _14779_/X sky130_fd_sc_hd__or2_1
XFILLER_32_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19306_ _19306_/CLK _19306_/D vssd1 vssd1 vccd1 vccd1 _19306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ _16551_/A0 _19124_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _19124_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17498_ _17498_/A _17547_/B vssd1 vssd1 vccd1 vccd1 _17498_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19237_ _19273_/CLK _19237_/D vssd1 vssd1 vccd1 vccd1 _19237_/Q sky130_fd_sc_hd__dfxtp_1
X_16449_ _19057_/Q _16614_/A0 _16454_/S vssd1 vssd1 vccd1 vccd1 _19057_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19168_ _19653_/A _19168_/D vssd1 vssd1 vccd1 vccd1 _19168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18119_ _18593_/CLK _18119_/D vssd1 vssd1 vccd1 vccd1 _18119_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_144_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19099_ _19099_/CLK _19099_/D vssd1 vssd1 vccd1 vccd1 _19099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09823_ _11691_/B1 _09991_/A _09822_/X _11692_/A1 _18375_/Q vssd1 vssd1 vccd1 vccd1
+ _09823_/X sky130_fd_sc_hd__o32a_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09754_ _11251_/S _19166_/Q _09770_/S _09753_/X vssd1 vssd1 vccd1 vccd1 _09754_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09685_ _09845_/S _09684_/X _10996_/B1 vssd1 vssd1 vccd1 vccd1 _09685_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10460_ _19643_/Q _18932_/Q _10613_/S vssd1 vssd1 vccd1 vccd1 _10460_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09119_ _19046_/Q _11167_/B _09919_/C1 _09118_/X vssd1 vssd1 vccd1 vccd1 _09119_/X
+ sky130_fd_sc_hd__a211o_1
X_10391_ _10866_/S _10389_/X _10390_/X vssd1 vssd1 vccd1 vccd1 _10391_/X sky130_fd_sc_hd__o21a_1
XFILLER_136_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ _17838_/Q _12130_/B vssd1 vssd1 vccd1 vccd1 _12136_/C sky130_fd_sc_hd__and2_2
XFILLER_124_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12061_ _17808_/Q _12085_/B vssd1 vssd1 vccd1 vccd1 _12061_/X sky130_fd_sc_hd__or2_1
Xfanout1903 _16110_/B1 vssd1 vssd1 vccd1 vccd1 _14991_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ _18829_/Q _11479_/B vssd1 vssd1 vccd1 vccd1 _11012_/X sky130_fd_sc_hd__or2_1
XFILLER_132_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15820_ _18612_/Q _17710_/A0 _15832_/S vssd1 vssd1 vccd1 vccd1 _18612_/D sky130_fd_sc_hd__mux2_1
Xfanout960 _14489_/Y vssd1 vssd1 vccd1 vccd1 _14521_/S sky130_fd_sc_hd__clkbuf_16
Xfanout971 _14070_/S vssd1 vssd1 vccd1 vccd1 _14072_/S sky130_fd_sc_hd__buf_12
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout982 _12762_/B vssd1 vssd1 vccd1 vccd1 _13579_/A sky130_fd_sc_hd__buf_6
XFILLER_77_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 _10531_/X vssd1 vssd1 vccd1 vccd1 _16418_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_253_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _15751_/A _15751_/B _15751_/C vssd1 vssd1 vccd1 vccd1 _15751_/X sky130_fd_sc_hd__or3_1
XFILLER_46_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12963_ _17827_/Q _13164_/A2 _13164_/B1 _17859_/Q vssd1 vssd1 vccd1 vccd1 _12963_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _12459_/X _13976_/B _14683_/X _18627_/Q vssd1 vssd1 vccd1 vccd1 _14702_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _19155_/CLK _18470_/D vssd1 vssd1 vccd1 vccd1 _18470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11914_ _18568_/Q _11918_/A2 _11706_/B _13081_/A vssd1 vssd1 vccd1 vccd1 _11914_/X
+ sky130_fd_sc_hd__a22o_4
X_15682_ _15744_/A _15725_/A vssd1 vssd1 vccd1 vccd1 _15684_/A sky130_fd_sc_hd__nor2_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12894_ _13134_/S _12811_/X _12746_/X vssd1 vssd1 vccd1 vccd1 _12895_/A sky130_fd_sc_hd__a21bo_1
XANTENNA_320 _18105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_331 _17124_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_342 _11482_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _18568_/Q _17461_/A2 _17426_/B1 vssd1 vssd1 vccd1 vccd1 _17421_/X sky130_fd_sc_hd__o21a_1
XFILLER_261_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14633_ _17692_/A0 _18439_/Q _14648_/S vssd1 vssd1 vccd1 vccd1 _18439_/D sky130_fd_sc_hd__mux2_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11845_ _11845_/A _11845_/B vssd1 vssd1 vccd1 vccd1 _11845_/X sky130_fd_sc_hd__or2_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 _09750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_364 _12320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_375 _14708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_386 _17208_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_397 _12599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _17352_/A _17352_/B vssd1 vssd1 vccd1 vccd1 _19473_/D sky130_fd_sc_hd__and2_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14592_/A _14564_/B vssd1 vssd1 vccd1 vccd1 _18390_/D sky130_fd_sc_hd__or2_1
XFILLER_220_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _12842_/A _12837_/B _11859_/A vssd1 vssd1 vccd1 vccd1 _11776_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_159_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _17701_/A0 _18916_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _18916_/D sky130_fd_sc_hd__mux2_1
XFILLER_202_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13515_ _13515_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13515_/Y sky130_fd_sc_hd__nor2_1
XFILLER_186_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17283_ _17498_/A _17250_/B _18122_/Q _17540_/B1 vssd1 vssd1 vccd1 vccd1 _17283_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10727_ _11618_/A1 _18226_/Q _10726_/S _18961_/Q _10745_/S vssd1 vssd1 vccd1 vccd1
+ _10727_/X sky130_fd_sc_hd__o221a_1
X_14495_ _17697_/A0 _18345_/Q _14517_/S vssd1 vssd1 vccd1 vccd1 _18345_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19022_ _19632_/CLK _19022_/D vssd1 vssd1 vccd1 vccd1 _19022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ _17698_/A0 _18849_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _18849_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13446_ _15450_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13446_/Y sky130_fd_sc_hd__nand2_1
X_10658_ _18259_/Q _18834_/Q _10667_/S vssd1 vssd1 vccd1 vccd1 _10658_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16165_ _17695_/A0 _18782_/Q _16165_/S vssd1 vssd1 vccd1 vccd1 _18782_/D sky130_fd_sc_hd__mux2_1
X_13377_ input269/X _12575_/Y _13371_/X _13427_/A1 vssd1 vssd1 vccd1 vccd1 _13377_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_155_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10589_ _10585_/X _10588_/X _10589_/S vssd1 vssd1 vccd1 vccd1 _10589_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15116_ _15116_/A _15116_/B _17556_/A vssd1 vssd1 vccd1 vccd1 _15123_/B sky130_fd_sc_hd__or3b_4
X_12328_ _17815_/Q _17814_/Q _17813_/Q _17812_/Q vssd1 vssd1 vccd1 vccd1 _12333_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_86_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16096_ _16096_/A1 _16095_/Y _16149_/A vssd1 vssd1 vccd1 vccd1 _18750_/D sky130_fd_sc_hd__a21oi_1
XFILLER_141_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15047_ _16459_/B _15047_/B vssd1 vssd1 vccd1 vccd1 _15047_/Y sky130_fd_sc_hd__nor2_8
X_12259_ _17886_/Q _12257_/B _12203_/A vssd1 vssd1 vccd1 vccd1 _12259_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_272_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18806_ _19623_/CLK _18806_/D vssd1 vssd1 vccd1 vccd1 _18806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16998_ _17573_/A _17044_/A2 _16997_/X _17559_/A vssd1 vssd1 vccd1 vccd1 _19335_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18737_ _18738_/CLK _18737_/D vssd1 vssd1 vccd1 vccd1 _18737_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_49_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15949_ _18692_/Q _15949_/A2 _15948_/X _14205_/A vssd1 vssd1 vccd1 vccd1 _18692_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09470_ _09350_/S _09467_/X _09460_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09470_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18668_ _18715_/CLK _18668_/D vssd1 vssd1 vccd1 vccd1 _18668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17619_ _19389_/Q _15092_/B input175/X _17592_/X _17623_/B1 vssd1 vssd1 vccd1 vccd1
+ _17619_/X sky130_fd_sc_hd__a41o_1
XFILLER_52_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18599_ _18880_/CLK _18599_/D vssd1 vssd1 vccd1 vccd1 _18599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19225_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09806_ _19070_/Q _18974_/Q _11617_/S vssd1 vssd1 vccd1 vccd1 _09806_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09737_ _11217_/A _09027_/A _09036_/X _09483_/Y _08999_/A vssd1 vssd1 vccd1 vccd1
+ _09737_/X sky130_fd_sc_hd__a32o_1
XFILLER_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09668_ _09666_/X _09667_/X _10315_/S vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__mux2_1
XFILLER_227_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09599_ _18053_/Q _10364_/B _09598_/X _09718_/S vssd1 vssd1 vccd1 vccd1 _09599_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _13908_/A _11555_/B _10160_/A vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__a21oi_4
XFILLER_202_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ _11566_/A1 _17789_/Q _11070_/S _18338_/Q vssd1 vssd1 vccd1 vccd1 _11561_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_156_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ _19436_/Q _12582_/X _13299_/X vssd1 vssd1 vccd1 vccd1 _13300_/X sky130_fd_sc_hd__o21a_1
X_10512_ _10662_/A1 _18158_/Q _18804_/Q _10582_/S vssd1 vssd1 vccd1 vccd1 _10512_/X
+ sky130_fd_sc_hd__a22o_1
X_14280_ _17698_/A0 _18139_/Q _14301_/S vssd1 vssd1 vccd1 vccd1 _18139_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11492_ _11513_/A1 _19598_/Q _19566_/Q _10424_/S vssd1 vssd1 vccd1 vccd1 _11492_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ _14156_/A0 _13230_/X _09230_/B vssd1 vssd1 vccd1 vccd1 _13231_/Y sky130_fd_sc_hd__o21ai_1
X_10443_ _10441_/X _10442_/X _10668_/S vssd1 vssd1 vccd1 vccd1 _10444_/B sky130_fd_sc_hd__mux2_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13162_ _15330_/A _13162_/B vssd1 vssd1 vccd1 vccd1 _13185_/C sky130_fd_sc_hd__nor2_1
XFILLER_163_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10374_ _10747_/A1 _10373_/X _08903_/A vssd1 vssd1 vccd1 vccd1 _10374_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12113_ _12203_/A _12113_/B _12114_/B vssd1 vssd1 vccd1 vccd1 _17831_/D sky130_fd_sc_hd__nor3_1
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17970_ _18627_/CLK _17970_/D vssd1 vssd1 vccd1 vccd1 _17970_/Q sky130_fd_sc_hd__dfxtp_1
X_13093_ _13414_/A _12817_/Y _12745_/X vssd1 vssd1 vccd1 vccd1 _13093_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1700 _09457_/A vssd1 vssd1 vccd1 vccd1 _09095_/A sky130_fd_sc_hd__buf_12
XFILLER_266_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16921_ _18761_/Q _16969_/A2 _16969_/B1 input225/X _16965_/C1 vssd1 vssd1 vccd1 vccd1
+ _16921_/X sky130_fd_sc_hd__a221o_2
X_12044_ _17897_/Q _12052_/A2 _12043_/X _13100_/A vssd1 vssd1 vccd1 vccd1 _17799_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1711 _08842_/Y vssd1 vssd1 vccd1 vccd1 _12488_/B sky130_fd_sc_hd__buf_12
XFILLER_78_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1722 _08825_/A vssd1 vssd1 vccd1 vccd1 _16020_/A sky130_fd_sc_hd__buf_4
Xfanout1733 _18658_/Q vssd1 vssd1 vccd1 vccd1 _15088_/B sky130_fd_sc_hd__clkbuf_4
Xfanout1744 _18273_/Q vssd1 vssd1 vccd1 vccd1 _15007_/S sky130_fd_sc_hd__buf_2
XFILLER_265_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19640_ _19640_/CLK _19640_/D vssd1 vssd1 vccd1 vccd1 _19640_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1755 _17912_/Q vssd1 vssd1 vccd1 vccd1 _11252_/S sky130_fd_sc_hd__buf_12
XFILLER_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16852_ _16852_/A _17922_/Q vssd1 vssd1 vccd1 vccd1 _16852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_277_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1766 _15129_/B2 vssd1 vssd1 vccd1 vccd1 _12466_/A0 sky130_fd_sc_hd__buf_12
XFILLER_226_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1777 _17908_/Q vssd1 vssd1 vccd1 vccd1 _09457_/B sky130_fd_sc_hd__buf_12
XFILLER_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout790 _16492_/Y vssd1 vssd1 vccd1 vccd1 _16515_/S sky130_fd_sc_hd__buf_6
Xfanout1788 _10513_/S vssd1 vssd1 vccd1 vccd1 _10036_/S sky130_fd_sc_hd__buf_6
X_15803_ _18595_/Q _17693_/A0 _15829_/S vssd1 vssd1 vccd1 vccd1 _18595_/D sky130_fd_sc_hd__mux2_1
Xfanout1799 _17804_/Q vssd1 vssd1 vccd1 vccd1 _12053_/A sky130_fd_sc_hd__buf_8
XFILLER_19_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16783_ _19282_/Q _19281_/Q _16783_/C vssd1 vssd1 vccd1 vccd1 _16786_/B sky130_fd_sc_hd__and3_1
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19571_ _19635_/CLK _19571_/D vssd1 vssd1 vccd1 vccd1 _19571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13995_ _14033_/A1 _13251_/X _13994_/X _16153_/D vssd1 vssd1 vccd1 vccd1 _17962_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18522_ _19286_/CLK _18522_/D vssd1 vssd1 vccd1 vccd1 _18522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15734_ _19484_/Q _19418_/Q vssd1 vssd1 vccd1 vccd1 _15757_/A sky130_fd_sc_hd__or2_1
XFILLER_46_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ _13135_/S _12941_/X _12945_/Y _13194_/S vssd1 vssd1 vccd1 vccd1 _12946_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ _19632_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_1
X_15665_ _15686_/B _15665_/B vssd1 vssd1 vccd1 vccd1 _15665_/X sky130_fd_sc_hd__xor2_1
XFILLER_222_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12877_ _12877_/A vssd1 vssd1 vccd1 vccd1 _12877_/Y sky130_fd_sc_hd__inv_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 _11868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_161 _12379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _13996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17404_ _17404_/A _17423_/B vssd1 vssd1 vccd1 vccd1 _17404_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _17708_/A0 _18423_/Q _14622_/S vssd1 vssd1 vccd1 vccd1 _18423_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_183 _14014_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ _11828_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11828_/X sky130_fd_sc_hd__or2_4
X_18384_ _19399_/CLK _18384_/D vssd1 vssd1 vccd1 vccd1 _18384_/Q sky130_fd_sc_hd__dfxtp_4
X_15596_ _18123_/Q _15763_/A2 _15595_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _15639_/B
+ sky130_fd_sc_hd__o22a_4
XANTENNA_194 _14028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _19465_/Q _17577_/A _17361_/S vssd1 vssd1 vccd1 vccd1 _17336_/B sky130_fd_sc_hd__mux2_1
XFILLER_186_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14547_ _18382_/Q _14575_/A2 _14575_/B1 input41/X vssd1 vssd1 vccd1 vccd1 _14548_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_230_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11759_ _18577_/Q _11759_/A2 _11844_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _11759_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17266_ _18116_/Q _17129_/A _17468_/A _17310_/B vssd1 vssd1 vccd1 vccd1 _17266_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14478_ _18330_/Q _17682_/A0 _14486_/S vssd1 vssd1 vccd1 vccd1 _18330_/D sky130_fd_sc_hd__mux2_1
X_16217_ _16614_/A0 _18833_/Q _16222_/S vssd1 vssd1 vccd1 vccd1 _18833_/D sky130_fd_sc_hd__mux2_1
X_19005_ _19133_/CLK _19005_/D vssd1 vssd1 vccd1 vccd1 _19005_/Q sky130_fd_sc_hd__dfxtp_1
X_13429_ _19505_/Q _13781_/A2 _13781_/B1 _13428_/X vssd1 vssd1 vccd1 vccd1 _13429_/X
+ sky130_fd_sc_hd__o211a_1
X_17197_ _19417_/Q fanout533/X _17517_/A _17119_/B vssd1 vssd1 vccd1 vccd1 _17198_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16148_ _14186_/S _16145_/C _16154_/A vssd1 vssd1 vccd1 vccd1 _16149_/B sky130_fd_sc_hd__o21a_1
XFILLER_143_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_171_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19453_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_100_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19157_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08970_ _09723_/S _08967_/X _08969_/X vssd1 vssd1 vccd1 vccd1 _08970_/Y sky130_fd_sc_hd__a21oi_4
X_16079_ _18742_/Q _16093_/B vssd1 vssd1 vccd1 vccd1 _16079_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 coreIndex[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_8
XFILLER_84_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09522_ _11622_/C1 _09516_/X _09519_/X _09521_/X _11495_/B1 vssd1 vssd1 vccd1 vccd1
+ _09523_/C sky130_fd_sc_hd__a311o_1
XFILLER_65_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09453_ _19625_/Q _18914_/Q _09464_/S vssd1 vssd1 vccd1 vccd1 _09453_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09384_ _18315_/Q _17766_/Q _10128_/B vssd1 vssd1 vccd1 vccd1 _09384_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput360 _11795_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[4] sky130_fd_sc_hd__buf_4
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput371 _08863_/Y vssd1 vssd1 vccd1 vccd1 core_wb_we_o sky130_fd_sc_hd__buf_4
XFILLER_105_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput382 _11935_/X vssd1 vssd1 vccd1 vccd1 din0[15] sky130_fd_sc_hd__buf_4
X_10090_ _18469_/Q _18370_/Q _10090_/S vssd1 vssd1 vccd1 vccd1 _10090_/X sky130_fd_sc_hd__mux2_1
Xfanout1007 _16485_/S vssd1 vssd1 vccd1 vccd1 _16491_/S sky130_fd_sc_hd__buf_8
Xoutput393 _11945_/X vssd1 vssd1 vccd1 vccd1 din0[25] sky130_fd_sc_hd__buf_4
XFILLER_121_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1018 _14384_/X vssd1 vssd1 vccd1 vccd1 _14402_/S sky130_fd_sc_hd__buf_12
Xfanout1029 _16530_/A0 vssd1 vssd1 vccd1 vccd1 _16431_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_259_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12800_ _12723_/X _12677_/X _12823_/A vssd1 vssd1 vccd1 vccd1 _12800_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13780_ _19548_/Q _13921_/S vssd1 vssd1 vccd1 vccd1 _13780_/X sky130_fd_sc_hd__or2_1
X_10992_ _18644_/Q _18066_/Q _11386_/S vssd1 vssd1 vccd1 vccd1 _10992_/X sky130_fd_sc_hd__mux2_1
XFILLER_262_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _12730_/Y _12728_/X _12821_/A vssd1 vssd1 vccd1 vccd1 _12731_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _15450_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _15450_/Y sky130_fd_sc_hd__nor2_1
XFILLER_203_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12662_ _13860_/B _12656_/X _12661_/X _11629_/B vssd1 vssd1 vccd1 vccd1 _12663_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14401_ _16542_/A0 _18252_/Q _14412_/S vssd1 vssd1 vccd1 vccd1 _18252_/D sky130_fd_sc_hd__mux2_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _18047_/Q _18015_/Q _11613_/S vssd1 vssd1 vccd1 vccd1 _11613_/X sky130_fd_sc_hd__mux2_1
X_15381_ _15404_/B _13363_/Y _15381_/A3 _15380_/X vssd1 vssd1 vccd1 vccd1 _15381_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_212_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12593_ _12593_/A _13568_/A vssd1 vssd1 vccd1 vccd1 _12593_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17120_ _17214_/A _17120_/B vssd1 vssd1 vccd1 vccd1 _17120_/Y sky130_fd_sc_hd__nand2_8
XFILLER_11_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14332_ _18189_/Q _17716_/A0 _14339_/S vssd1 vssd1 vccd1 vccd1 _18189_/D sky130_fd_sc_hd__mux2_1
X_11544_ _11545_/B _10603_/A _11545_/A vssd1 vssd1 vccd1 vccd1 _11544_/X sky130_fd_sc_hd__o21ba_1
XFILLER_184_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ _17051_/A _17051_/B _17051_/C _17051_/D vssd1 vssd1 vccd1 vccd1 _17052_/D
+ sky130_fd_sc_hd__or4_1
X_14263_ _18303_/Q _14267_/A2 _14262_/X _14451_/B vssd1 vssd1 vccd1 vccd1 _18129_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11475_ _12488_/B _11468_/Y _11470_/Y _11474_/Y _08843_/Y vssd1 vssd1 vccd1 vccd1
+ _11475_/X sky130_fd_sc_hd__a311o_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16002_ _18716_/Q _16002_/A2 _16002_/B1 _18765_/Q _16002_/C1 vssd1 vssd1 vccd1 vccd1
+ _16002_/X sky130_fd_sc_hd__a221o_1
X_13214_ _15884_/A _12506_/X _13206_/X _13213_/X _12510_/X vssd1 vssd1 vccd1 vccd1
+ _13214_/X sky130_fd_sc_hd__o221a_1
XFILLER_7_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10426_ _19093_/Q _18997_/Q _10426_/S vssd1 vssd1 vccd1 vccd1 _10426_/X sky130_fd_sc_hd__mux2_1
X_14194_ _18708_/Q _18095_/Q _14200_/S vssd1 vssd1 vccd1 vccd1 _14195_/B sky130_fd_sc_hd__mux2_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13145_ _09405_/Y _13292_/A2 _13144_/X _13256_/B1 _17927_/Q vssd1 vssd1 vccd1 vccd1
+ _13146_/B sky130_fd_sc_hd__a32o_1
X_10357_ _11046_/S1 _10346_/X _10356_/X _11438_/B1 vssd1 vssd1 vccd1 vccd1 _10357_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _17982_/CLK _17953_/D vssd1 vssd1 vccd1 vccd1 _17953_/Q sky130_fd_sc_hd__dfxtp_1
X_13076_ _13986_/B vssd1 vssd1 vccd1 vccd1 _13076_/Y sky130_fd_sc_hd__inv_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10288_ _10294_/A1 _19223_/Q _19191_/Q _10299_/S _10293_/B1 vssd1 vssd1 vccd1 vccd1
+ _10288_/X sky130_fd_sc_hd__a221o_1
XFILLER_266_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16904_ _16904_/A _16904_/B vssd1 vssd1 vccd1 vccd1 _19310_/D sky130_fd_sc_hd__and2_1
X_12027_ _17791_/Q _12051_/B vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__or2_1
Xfanout1530 _11189_/A vssd1 vssd1 vccd1 vccd1 _11282_/A sky130_fd_sc_hd__buf_6
XFILLER_239_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1541 _08900_/Y vssd1 vssd1 vccd1 vccd1 _10653_/A1 sky130_fd_sc_hd__buf_12
X_17884_ _19261_/CLK _17884_/D vssd1 vssd1 vccd1 vccd1 _17884_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1552 _10280_/S vssd1 vssd1 vccd1 vccd1 _09723_/S sky130_fd_sc_hd__buf_8
XFILLER_120_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1563 _11515_/B1 vssd1 vssd1 vccd1 vccd1 _08903_/A sky130_fd_sc_hd__buf_8
Xfanout1574 _11198_/S vssd1 vssd1 vccd1 vccd1 _11285_/S sky130_fd_sc_hd__buf_8
XFILLER_239_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19623_ _19623_/CLK _19623_/D vssd1 vssd1 vccd1 vccd1 _19623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16835_ _17814_/Q _14682_/A _16836_/S vssd1 vssd1 vccd1 vccd1 _17051_/D sky130_fd_sc_hd__mux2_1
Xfanout1585 _11274_/S1 vssd1 vssd1 vccd1 vccd1 _11622_/A1 sky130_fd_sc_hd__buf_6
Xfanout1596 _08894_/Y vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__buf_12
XFILLER_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19554_ _19586_/CLK _19554_/D vssd1 vssd1 vccd1 vccd1 _19554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16766_ _19275_/Q _16767_/C _19276_/Q vssd1 vssd1 vccd1 vccd1 _16768_/B sky130_fd_sc_hd__a21oi_1
X_13978_ _14004_/A _13978_/B vssd1 vssd1 vccd1 vccd1 _13978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18505_ _19229_/CLK _18505_/D vssd1 vssd1 vccd1 vccd1 _18505_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15717_ _15709_/X _15710_/X _15716_/X _15717_/B2 _15782_/B1 vssd1 vssd1 vccd1 vccd1
+ _15717_/X sky130_fd_sc_hd__a221o_1
X_12929_ _13079_/A _12923_/Y _12924_/X _12928_/X vssd1 vssd1 vccd1 vccd1 _12929_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_280_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16697_ _19252_/Q _16697_/B vssd1 vssd1 vccd1 vccd1 _16704_/C sky130_fd_sc_hd__and2_1
X_19485_ _19485_/CLK _19485_/D vssd1 vssd1 vccd1 vccd1 _19485_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18436_ _19615_/CLK _18436_/D vssd1 vssd1 vccd1 vccd1 _18436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15648_ _15623_/A _15645_/X _15647_/X vssd1 vssd1 vccd1 vccd1 _15648_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18367_ _19645_/CLK _18367_/D vssd1 vssd1 vccd1 vccd1 _18367_/Q sky130_fd_sc_hd__dfxtp_1
X_15579_ _15580_/A _15580_/B _15638_/B vssd1 vssd1 vccd1 vccd1 _15579_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_187_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17318_ _17378_/A _17318_/B vssd1 vssd1 vccd1 vccd1 _19456_/D sky130_fd_sc_hd__and2_1
XFILLER_179_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18298_ _19444_/CLK _18298_/D vssd1 vssd1 vccd1 vccd1 _18298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17249_ _17247_/Y _17248_/X _17261_/A vssd1 vssd1 vccd1 vccd1 _19433_/D sky130_fd_sc_hd__a21oi_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08953_ _08903_/A _14488_/C _14074_/C _09498_/S _08956_/B vssd1 vssd1 vccd1 vccd1
+ _08954_/C sky130_fd_sc_hd__o221a_1
XFILLER_229_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08884_ _18406_/Q _18405_/Q vssd1 vssd1 vccd1 vccd1 _08884_/X sky130_fd_sc_hd__or2_4
XFILLER_257_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ _12389_/A1 _09492_/X _09493_/X vssd1 vssd1 vccd1 vccd1 _09505_/X sky130_fd_sc_hd__o21a_1
XFILLER_225_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09866_/B _15238_/A _09405_/Y vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__o21a_4
XFILLER_213_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09367_ _18109_/Q _09367_/B vssd1 vssd1 vccd1 vccd1 _09367_/X sky130_fd_sc_hd__or2_2
XFILLER_178_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09298_ _18316_/Q _17767_/Q _09306_/S vssd1 vssd1 vccd1 vccd1 _09298_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_50 _12613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_61 _10121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_83 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_94 _10913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11260_ _12595_/A vssd1 vssd1 vccd1 vccd1 _11292_/A sky130_fd_sc_hd__inv_2
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10211_ _10211_/A1 _10205_/X _10208_/X _11053_/A vssd1 vssd1 vccd1 vccd1 _10211_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_137_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191_ _08901_/A _19115_/Q _19147_/Q _09883_/B vssd1 vssd1 vccd1 vccd1 _11191_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10142_ _10140_/X _10141_/X _10225_/S vssd1 vssd1 vccd1 vccd1 _10142_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ _14946_/Y _14949_/X _14950_/B1 vssd1 vssd1 vccd1 vccd1 _14950_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10073_ _11739_/A _11739_/B _09560_/X _13044_/S vssd1 vssd1 vccd1 vccd1 _10074_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13901_ _18129_/Q _13900_/C _18130_/Q vssd1 vssd1 vccd1 vccd1 _13902_/B sky130_fd_sc_hd__a21oi_1
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14881_ _15003_/A1 _13561_/Y _15003_/B1 _18645_/Q _15003_/C1 vssd1 vssd1 vccd1 vccd1
+ _14881_/X sky130_fd_sc_hd__a221o_1
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16620_ _17720_/A0 _19223_/Q _16622_/S vssd1 vssd1 vccd1 vccd1 _19223_/D sky130_fd_sc_hd__mux2_1
X_13832_ _13637_/A _14028_/B _13818_/X vssd1 vssd1 vccd1 vccd1 _13832_/X sky130_fd_sc_hd__o21a_1
XFILLER_223_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16551_ _16551_/A0 _19156_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _19156_/D sky130_fd_sc_hd__mux2_1
XFILLER_216_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13763_ _13763_/A _13763_/B vssd1 vssd1 vccd1 vccd1 _14150_/A sky130_fd_sc_hd__xnor2_2
XFILLER_44_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10975_ _11358_/A _10970_/X _10974_/X vssd1 vssd1 vccd1 vccd1 _10977_/C sky130_fd_sc_hd__a21oi_1
XFILLER_204_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12714_ _12612_/B _12650_/B _12733_/S vssd1 vssd1 vccd1 vccd1 _12714_/X sky130_fd_sc_hd__mux2_1
X_15502_ _15502_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _15502_/Y sky130_fd_sc_hd__nor2_1
XFILLER_280_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19270_ _19273_/CLK _19270_/D vssd1 vssd1 vccd1 vccd1 _19270_/Q sky130_fd_sc_hd__dfxtp_1
X_16482_ _16548_/A0 _19089_/Q _16485_/S vssd1 vssd1 vccd1 vccd1 _19089_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13694_ _13931_/A _13692_/Y _13693_/X _13695_/A _13294_/A vssd1 vssd1 vccd1 vccd1
+ _13694_/X sky130_fd_sc_hd__o32a_1
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15433_ _15456_/C _15410_/B _15407_/X vssd1 vssd1 vccd1 vccd1 _15436_/B sky130_fd_sc_hd__o21ai_1
X_18221_ _19118_/CLK _18221_/D vssd1 vssd1 vccd1 vccd1 _18221_/Q sky130_fd_sc_hd__dfxtp_1
X_12645_ _10677_/A _10675_/Y _12644_/Y vssd1 vssd1 vccd1 vccd1 _12645_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18152_ _19632_/CLK _18152_/D vssd1 vssd1 vccd1 vccd1 _18152_/Q sky130_fd_sc_hd__dfxtp_1
X_15364_ _15364_/A _15364_/B vssd1 vssd1 vccd1 vccd1 _15364_/Y sky130_fd_sc_hd__nand2_1
X_12576_ _12576_/A _12576_/B vssd1 vssd1 vccd1 vccd1 _12859_/S sky130_fd_sc_hd__or2_4
XFILLER_200_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14315_ _18172_/Q _16500_/A0 _14335_/S vssd1 vssd1 vccd1 vccd1 _18172_/D sky130_fd_sc_hd__mux2_1
X_17103_ _19385_/Q _17115_/B vssd1 vssd1 vccd1 vccd1 _17103_/X sky130_fd_sc_hd__or2_1
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18083_ _19304_/CLK _18083_/D vssd1 vssd1 vccd1 vccd1 _18083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11527_ _13351_/A _11680_/B _13357_/S vssd1 vssd1 vccd1 vccd1 _11679_/B sky130_fd_sc_hd__a21oi_4
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15295_ _15307_/B _15292_/X _15294_/Y _15416_/A vssd1 vssd1 vccd1 vccd1 _15295_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17034_ _17196_/B _17046_/A2 _17033_/X _17106_/C1 vssd1 vssd1 vccd1 vccd1 _19353_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14246_ _18121_/Q _14266_/B vssd1 vssd1 vccd1 vccd1 _14246_/X sky130_fd_sc_hd__or2_1
XFILLER_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11458_ _11458_/A1 _19143_/Q _11462_/S _19111_/Q _10403_/S vssd1 vssd1 vccd1 vccd1
+ _11458_/X sky130_fd_sc_hd__o221a_1
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10409_ _10409_/A _10409_/B vssd1 vssd1 vccd1 vccd1 _10409_/X sky130_fd_sc_hd__or2_2
XFILLER_194_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14177_ _14177_/A _14177_/B vssd1 vssd1 vccd1 vccd1 _18086_/D sky130_fd_sc_hd__and2_1
X_11389_ _11389_/A1 _17771_/Q _11386_/S _18320_/Q _10403_/S vssd1 vssd1 vccd1 vccd1
+ _11389_/X sky130_fd_sc_hd__o221a_1
XFILLER_259_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13224_/B _14143_/A _13125_/X _12442_/C vssd1 vssd1 vccd1 vccd1 _13128_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_12__f_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_91_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _19118_/CLK _18985_/D vssd1 vssd1 vccd1 vccd1 _18985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13059_ _17829_/Q _13164_/A2 _13164_/B1 _17861_/Q vssd1 vssd1 vccd1 vccd1 _13059_/X
+ sky130_fd_sc_hd__a22o_1
X_17936_ _18660_/CLK _17936_/D vssd1 vssd1 vccd1 vccd1 _17936_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1360 _10101_/B vssd1 vssd1 vccd1 vccd1 _11479_/B sky130_fd_sc_hd__buf_6
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1371 _09843_/S vssd1 vssd1 vccd1 vccd1 _10856_/C sky130_fd_sc_hd__buf_4
X_17867_ _19300_/CLK _17867_/D vssd1 vssd1 vccd1 vccd1 _17867_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1382 fanout1386/X vssd1 vssd1 vccd1 vccd1 _11247_/S sky130_fd_sc_hd__buf_6
Xfanout1393 _10320_/S vssd1 vssd1 vccd1 vccd1 _11171_/S sky130_fd_sc_hd__buf_6
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19606_ _19649_/CLK _19606_/D vssd1 vssd1 vccd1 vccd1 _19606_/Q sky130_fd_sc_hd__dfxtp_1
X_16818_ _08821_/Y _16816_/C _16817_/Y vssd1 vssd1 vccd1 vccd1 _19295_/D sky130_fd_sc_hd__a21oi_1
X_17798_ _18201_/CLK _17798_/D vssd1 vssd1 vccd1 vccd1 _17798_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_207_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19537_ _19537_/CLK _19537_/D vssd1 vssd1 vccd1 vccd1 _19537_/Q sky130_fd_sc_hd__dfxtp_1
X_16749_ _19269_/Q _16751_/C _16748_/Y vssd1 vssd1 vccd1 vccd1 _19269_/D sky130_fd_sc_hd__a21oi_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19468_ _19502_/CLK _19468_/D vssd1 vssd1 vccd1 vccd1 _19468_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_250_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09221_ _10200_/S _09214_/X _09213_/X _10356_/C1 vssd1 vssd1 vccd1 vccd1 _09221_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_222_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18419_ _19630_/CLK _18419_/D vssd1 vssd1 vccd1 vccd1 _18419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19399_ _19399_/CLK _19399_/D vssd1 vssd1 vccd1 vccd1 _19399_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_148_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09152_ _09027_/A _10085_/B _09148_/X _09151_/X _09019_/Y vssd1 vssd1 vccd1 vccd1
+ _09152_/X sky130_fd_sc_hd__a32o_1
XFILLER_148_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09083_ _09083_/A _13916_/A vssd1 vssd1 vccd1 vccd1 _15082_/B sky130_fd_sc_hd__nand2_8
XFILLER_238_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput70 dout0[34] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_2
XFILLER_238_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput81 dout0[44] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput92 dout0[54] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09985_ _17952_/Q _11295_/A2 _11216_/B1 vssd1 vssd1 vccd1 vccd1 _09985_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_104_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08936_ _08933_/X _08935_/X _08942_/B _08914_/X vssd1 vssd1 vccd1 vccd1 _08939_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08867_ _17891_/Q _17890_/Q _12267_/A vssd1 vssd1 vccd1 vccd1 _12443_/A sky130_fd_sc_hd__or3_4
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_wb_clk_i _19652_/A vssd1 vssd1 vccd1 vccd1 _19635_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10760_ _17941_/Q _08948_/B _10759_/X _08947_/B vssd1 vssd1 vccd1 vccd1 _10760_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09419_ _09718_/S _09419_/B vssd1 vssd1 vccd1 vccd1 _09424_/A sky130_fd_sc_hd__and2_1
XFILLER_158_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10691_ _18616_/Q _18187_/Q _11249_/S vssd1 vssd1 vccd1 vccd1 _10691_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12430_ _12430_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _12430_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12361_ _12420_/A1 _09991_/A _09012_/C _12420_/B1 _18380_/Q vssd1 vssd1 vccd1 vccd1
+ _12361_/X sky130_fd_sc_hd__o32a_1
XFILLER_139_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14100_ _17683_/A0 _18040_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _18040_/D sky130_fd_sc_hd__mux2_1
X_11312_ _11312_/A1 _17772_/Q _10940_/S _18321_/Q _10784_/S vssd1 vssd1 vccd1 vccd1
+ _11312_/X sky130_fd_sc_hd__o221a_1
X_15080_ _15081_/A _15120_/B vssd1 vssd1 vccd1 vccd1 _15080_/Y sky130_fd_sc_hd__nor2_1
X_12292_ _14681_/C _14682_/A _12292_/C vssd1 vssd1 vccd1 vccd1 _14688_/B sky130_fd_sc_hd__or3_2
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14031_ _17980_/Q _14032_/B _14030_/Y _16153_/D vssd1 vssd1 vccd1 vccd1 _17980_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11243_ _11251_/S _11250_/A1 _19210_/Q _09750_/S vssd1 vssd1 vccd1 vccd1 _11243_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11174_ _11168_/X _11170_/X _11173_/X _11406_/B2 _09350_/S vssd1 vssd1 vccd1 vccd1
+ _11174_/X sky130_fd_sc_hd__o221a_1
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10125_ _10123_/X _10124_/X _10200_/S vssd1 vssd1 vccd1 vccd1 _10125_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18770_ _18772_/CLK _18770_/D vssd1 vssd1 vccd1 vccd1 _18770_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15982_ _18706_/Q _16016_/A2 _16147_/A2 _18755_/Q _16018_/C1 vssd1 vssd1 vccd1 vccd1
+ _15982_/X sky130_fd_sc_hd__a221o_1
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17721_ _17721_/A0 _19647_/Q _17722_/S vssd1 vssd1 vccd1 vccd1 _19647_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10056_ _11282_/A _10054_/X _10055_/X _11285_/S vssd1 vssd1 vccd1 vccd1 _10056_/X
+ sky130_fd_sc_hd__a211o_1
X_14933_ _14931_/X _14932_/X _14714_/B vssd1 vssd1 vccd1 vccd1 _14933_/X sky130_fd_sc_hd__a21o_1
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _17685_/A0 _19580_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _19580_/D sky130_fd_sc_hd__mux2_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14864_ _18118_/Q _14893_/S _14852_/X _14863_/X vssd1 vssd1 vccd1 vccd1 _14864_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _09105_/A _19206_/Q _16622_/S vssd1 vssd1 vccd1 vccd1 _19206_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13815_ _13812_/A _12265_/B _13814_/X vssd1 vssd1 vccd1 vccd1 _13815_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_263_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17583_ _17583_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17583_/X sky130_fd_sc_hd__or2_1
X_14795_ _14795_/A vssd1 vssd1 vccd1 vccd1 _14795_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19322_ _19323_/CLK _19322_/D vssd1 vssd1 vccd1 vccd1 _19322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16534_ _17667_/A0 _19139_/Q _16556_/S vssd1 vssd1 vccd1 vccd1 _19139_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13746_ _17848_/Q _13821_/B vssd1 vssd1 vccd1 vccd1 _13746_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10958_ _11611_/S _10958_/B vssd1 vssd1 vccd1 vccd1 _10963_/A sky130_fd_sc_hd__and2_1
XFILLER_188_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19253_ _19261_/CLK _19253_/D vssd1 vssd1 vccd1 vccd1 _19253_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_204_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16465_ _16465_/A0 _19072_/Q _16485_/S vssd1 vssd1 vccd1 vccd1 _19072_/D sky130_fd_sc_hd__mux2_1
X_13677_ _12320_/A _13971_/A2 _13675_/Y _13676_/Y _13579_/A vssd1 vssd1 vccd1 vccd1
+ _13677_/X sky130_fd_sc_hd__a221o_4
X_10889_ _11596_/A1 _18153_/Q _18799_/Q _10815_/B vssd1 vssd1 vccd1 vccd1 _10889_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18204_ _19099_/CLK _18204_/D vssd1 vssd1 vccd1 vccd1 _18204_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12628_ _13357_/S _11446_/B _12625_/Y vssd1 vssd1 vccd1 vccd1 _12628_/X sky130_fd_sc_hd__o21a_1
X_15416_ _15416_/A _15416_/B _15416_/C vssd1 vssd1 vccd1 vccd1 _15416_/X sky130_fd_sc_hd__or3_1
X_19184_ _19216_/CLK _19184_/D vssd1 vssd1 vccd1 vccd1 _19184_/Q sky130_fd_sc_hd__dfxtp_1
X_16396_ _16594_/A0 _19005_/Q _16425_/S vssd1 vssd1 vccd1 vccd1 _19005_/D sky130_fd_sc_hd__mux2_1
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18135_ _19133_/CLK _18135_/D vssd1 vssd1 vccd1 vccd1 _18135_/Q sky130_fd_sc_hd__dfxtp_1
X_15347_ _15347_/A _15347_/B vssd1 vssd1 vccd1 vccd1 _15347_/Y sky130_fd_sc_hd__xnor2_1
X_12559_ _13167_/A _12561_/B vssd1 vssd1 vccd1 vccd1 _12559_/X sky130_fd_sc_hd__or2_1
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18066_ _19599_/CLK _18066_/D vssd1 vssd1 vccd1 vccd1 _18066_/Q sky130_fd_sc_hd__dfxtp_1
X_15278_ _19463_/Q _19397_/Q _15254_/B vssd1 vssd1 vccd1 vccd1 _15278_/X sky130_fd_sc_hd__a21o_1
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14229_ _18286_/Q _14247_/A2 _14228_/X _14450_/B vssd1 vssd1 vccd1 vccd1 _18112_/D
+ sky130_fd_sc_hd__o211a_1
X_17017_ _19345_/Q _17045_/B vssd1 vssd1 vccd1 vccd1 _17017_/X sky130_fd_sc_hd__or2_1
XFILLER_217_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_78_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19047_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout608 _13247_/C1 vssd1 vssd1 vccd1 vccd1 _13951_/C1 sky130_fd_sc_hd__buf_8
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout619 _17158_/B2 vssd1 vssd1 vccd1 vccd1 _17120_/B sky130_fd_sc_hd__buf_6
XFILLER_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09770_ _19621_/Q _18910_/Q _09770_/S vssd1 vssd1 vccd1 vccd1 _09770_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18968_ _19613_/CLK _18968_/D vssd1 vssd1 vccd1 vccd1 _18968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_258_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17919_ _18817_/CLK _17919_/D vssd1 vssd1 vccd1 vccd1 _17919_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18899_ _19219_/CLK _18899_/D vssd1 vssd1 vccd1 vccd1 _18899_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1190 _16002_/B1 vssd1 vssd1 vccd1 vccd1 _15976_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09204_ _09708_/A _09201_/X _09203_/Y _08895_/A vssd1 vssd1 vccd1 vccd1 _09204_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09135_ _09131_/X _09134_/X _09135_/S vssd1 vssd1 vccd1 vccd1 _09135_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09066_ _17901_/Q _12442_/B _11647_/A vssd1 vssd1 vccd1 vccd1 _09080_/B sky130_fd_sc_hd__and3_4
XFILLER_108_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09968_ _11190_/A1 _19555_/Q _09973_/S _19587_/Q _09972_/S vssd1 vssd1 vccd1 vccd1
+ _09968_/X sky130_fd_sc_hd__o221a_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ _08816_/A _17800_/Q vssd1 vssd1 vccd1 vccd1 _14306_/C sky130_fd_sc_hd__nand2b_2
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ _08939_/A _08939_/B _08939_/C _09042_/A _09042_/B vssd1 vssd1 vccd1 vccd1
+ _09899_/X sky130_fd_sc_hd__a32o_4
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _11810_/A _11944_/A1 _11814_/C _11959_/A2 input216/X vssd1 vssd1 vccd1 vccd1
+ _11930_/X sky130_fd_sc_hd__a32o_4
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_502 _15129_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_513 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ _11859_/A _11896_/A _11826_/A vssd1 vssd1 vccd1 vccd1 _11861_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_524 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_535 input220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13600_ _13797_/A0 _12756_/Y _13600_/S vssd1 vssd1 vccd1 vccd1 _13600_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_546 _15481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10812_ _19056_/Q _19024_/Q _10815_/B vssd1 vssd1 vccd1 vccd1 _10812_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14592_/A _14580_/B vssd1 vssd1 vccd1 vccd1 _18398_/D sky130_fd_sc_hd__or2_1
X_11792_ _11799_/A _11799_/B wire989/X vssd1 vssd1 vccd1 vccd1 _11792_/X sky130_fd_sc_hd__and3_1
XFILLER_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ _13545_/B _13961_/A vssd1 vssd1 vccd1 vccd1 _13531_/Y sky130_fd_sc_hd__nand2_1
X_10743_ _18461_/Q _18362_/Q _10744_/S vssd1 vssd1 vccd1 vccd1 _10743_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ _17714_/A0 _18865_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _18865_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _13462_/A _13462_/B _13462_/C vssd1 vssd1 vccd1 vccd1 _13462_/X sky130_fd_sc_hd__and3_2
X_10674_ _14252_/A _13679_/A _13739_/A vssd1 vssd1 vccd1 vccd1 _12729_/A sky130_fd_sc_hd__mux2_8
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15201_ _15199_/A _15199_/B _15200_/A vssd1 vssd1 vccd1 vccd1 _15201_/X sky130_fd_sc_hd__a21o_1
X_12413_ _10243_/A _12412_/A _12412_/Y _14001_/C1 vssd1 vssd1 vccd1 vccd1 _17912_/D
+ sky130_fd_sc_hd__o211a_1
X_16181_ _16611_/A0 _18798_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _18798_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13393_ _13387_/A _14155_/B _13392_/Y _11369_/B vssd1 vssd1 vccd1 vccd1 _13393_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_126_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15132_ _15133_/A _15133_/B vssd1 vssd1 vccd1 vccd1 _15132_/X sky130_fd_sc_hd__and2_4
X_12344_ _17889_/Q _12382_/A _12343_/Y _12350_/C1 vssd1 vssd1 vccd1 vccd1 _17889_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15063_ _18547_/Q _17707_/A0 _15070_/S vssd1 vssd1 vccd1 vccd1 _18547_/D sky130_fd_sc_hd__mux2_1
X_12275_ _16143_/C _16093_/B vssd1 vssd1 vccd1 vccd1 _12276_/B sky130_fd_sc_hd__nor2_4
XFILLER_175_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14014_ _14020_/B _14014_/B vssd1 vssd1 vccd1 vccd1 _14014_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11226_ _18641_/Q _18063_/Q _11226_/S vssd1 vssd1 vccd1 vccd1 _11226_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18822_ _18884_/CLK _18822_/D vssd1 vssd1 vccd1 vccd1 _18822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11157_ _11157_/A1 _17774_/Q _11154_/S _18323_/Q _10706_/S vssd1 vssd1 vccd1 vccd1
+ _11157_/X sky130_fd_sc_hd__o221a_1
XFILLER_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10108_ _10334_/A1 _17788_/Q _10090_/S _18337_/Q vssd1 vssd1 vccd1 vccd1 _10108_/X
+ sky130_fd_sc_hd__o22a_1
X_18753_ _18776_/CLK _18753_/D vssd1 vssd1 vccd1 vccd1 _18753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15965_ _18698_/Q _15977_/A2 _15964_/X _16968_/A vssd1 vssd1 vccd1 vccd1 _18698_/D
+ sky130_fd_sc_hd__o211a_1
X_11088_ _09457_/A _11085_/X _11087_/X vssd1 vssd1 vccd1 vccd1 _11088_/X sky130_fd_sc_hd__a21o_1
Xinput260 manufacturerID[6] vssd1 vssd1 vccd1 vccd1 _15875_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput271 partID[1] vssd1 vssd1 vccd1 vccd1 _15893_/A sky130_fd_sc_hd__clkbuf_2
X_17704_ _17704_/A0 _19630_/Q _17722_/S vssd1 vssd1 vccd1 vccd1 _19630_/D sky130_fd_sc_hd__mux2_1
Xinput282 versionID[2] vssd1 vssd1 vccd1 vccd1 _12851_/A sky130_fd_sc_hd__buf_2
XFILLER_264_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14916_ input57/X input92/X _14947_/S vssd1 vssd1 vccd1 vccd1 _14917_/A sky130_fd_sc_hd__mux2_2
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10039_ _19618_/Q _18907_/Q _11613_/S vssd1 vssd1 vccd1 vccd1 _10039_/X sky130_fd_sc_hd__mux2_1
X_18684_ _18691_/CLK _18684_/D vssd1 vssd1 vccd1 vccd1 _18684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_196_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19638_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15896_ input272/X _15941_/S vssd1 vssd1 vccd1 vccd1 _15896_/Y sky130_fd_sc_hd__nand2b_1
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17635_ _17668_/A0 _19563_/Q _17654_/S vssd1 vssd1 vccd1 vccd1 _19563_/D sky130_fd_sc_hd__mux2_1
XFILLER_223_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_125_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19321_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14847_ _14843_/Y _14846_/X _14879_/B1 vssd1 vssd1 vccd1 vccd1 _14847_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17566_ _19525_/Q _17561_/B _17588_/B1 _17565_/Y vssd1 vssd1 vccd1 vccd1 _19525_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14778_ _18479_/Q _14889_/B1 _14777_/Y _12243_/A vssd1 vssd1 vccd1 vccd1 _18479_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_223_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19305_ _19306_/CLK _19305_/D vssd1 vssd1 vccd1 vccd1 _19305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16517_ _10532_/B _19123_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _19123_/D sky130_fd_sc_hd__mux2_1
X_13729_ _13740_/B _13761_/B _13728_/Y vssd1 vssd1 vccd1 vccd1 _13729_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17497_ _18122_/Q _17539_/C1 _17495_/X _17496_/X vssd1 vssd1 vccd1 vccd1 _17497_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19236_ _19273_/CLK _19236_/D vssd1 vssd1 vccd1 vccd1 _19236_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16448_ _19056_/Q _16580_/A0 _16453_/S vssd1 vssd1 vccd1 vccd1 _19056_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19167_ _19622_/CLK _19167_/D vssd1 vssd1 vccd1 vccd1 _19167_/Q sky130_fd_sc_hd__dfxtp_1
X_16379_ _17711_/A0 _18990_/Q _16391_/S vssd1 vssd1 vccd1 vccd1 _18990_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18118_ _18593_/CLK _18118_/D vssd1 vssd1 vccd1 vccd1 _18118_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19098_ _19163_/CLK _19098_/D vssd1 vssd1 vccd1 vccd1 _19098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18049_ _19587_/CLK _18049_/D vssd1 vssd1 vccd1 vccd1 _18049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09822_ input129/X input134/X _09990_/S vssd1 vssd1 vccd1 vccd1 _09822_/X sky130_fd_sc_hd__mux2_8
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09753_ _11251_/S _11565_/A1 _19198_/Q _09750_/S vssd1 vssd1 vccd1 vccd1 _09753_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_274_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09684_ _18630_/Q _18052_/Q _19071_/Q _18975_/Q _11160_/S _10337_/S1 vssd1 vssd1
+ vccd1 vccd1 _09684_/X sky130_fd_sc_hd__mux4_1
XFILLER_255_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ _09457_/B _19014_/Q _09285_/C vssd1 vssd1 vccd1 vccd1 _09118_/X sky130_fd_sc_hd__and3_1
XFILLER_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10390_ _11312_/A1 _19221_/Q _19189_/Q _10864_/S _11584_/C1 vssd1 vssd1 vccd1 vccd1
+ _10390_/X sky130_fd_sc_hd__a221o_1
XFILLER_136_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09049_ _11141_/A _09050_/B vssd1 vssd1 vccd1 vccd1 _09049_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12060_ _08874_/D _12086_/A2 _12059_/X _14340_/A vssd1 vssd1 vccd1 vccd1 _17807_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11011_ _10243_/A _11006_/X _11010_/X _12466_/A0 vssd1 vssd1 vccd1 vccd1 _11011_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout1904 fanout1905/X vssd1 vssd1 vccd1 vccd1 _16110_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout950 _14660_/S vssd1 vssd1 vccd1 vccd1 _14663_/S sky130_fd_sc_hd__buf_12
XFILLER_77_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout961 _14108_/Y vssd1 vssd1 vccd1 vccd1 _14140_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout972 _14041_/Y vssd1 vssd1 vccd1 vccd1 _14070_/S sky130_fd_sc_hd__buf_12
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout983 _13808_/C1 vssd1 vssd1 vccd1 vccd1 _12762_/B sky130_fd_sc_hd__buf_8
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 _10531_/X vssd1 vssd1 vccd1 vccd1 _17683_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _15789_/A1 _15749_/Y _15789_/B1 vssd1 vssd1 vccd1 vccd1 _15751_/C sky130_fd_sc_hd__a21oi_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12962_ _12962_/A0 _15173_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _12962_/X sky130_fd_sc_hd__mux2_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _18471_/Q _14720_/A _14700_/Y _17159_/A vssd1 vssd1 vccd1 vccd1 _18471_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11913_ _18567_/Q _11918_/A2 _11706_/B _11740_/Y vssd1 vssd1 vccd1 vccd1 _11913_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_261_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_310 _18113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _18127_/Q _15763_/A2 _15680_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _15725_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12893_ _09897_/Y _13230_/A1 _12892_/Y _11731_/B vssd1 vssd1 vccd1 vccd1 _12899_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 _18105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_332 _11810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _13081_/A _17445_/A2 _17445_/B1 _17796_/Q _15116_/B vssd1 vssd1 vccd1 vccd1
+ _17420_/X sky130_fd_sc_hd__a221o_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _16426_/A _17691_/B vssd1 vssd1 vccd1 vccd1 _14632_/Y sky130_fd_sc_hd__nand2_2
XANTENNA_343 _11300_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ _11844_/A _11844_/B vssd1 vssd1 vccd1 vccd1 _11844_/X sky130_fd_sc_hd__and2_1
XFILLER_260_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_354 _12488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_365 _10373_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_376 _14807_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_387 _17208_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _19473_/Q _17172_/B _17361_/S vssd1 vssd1 vccd1 vccd1 _17352_/B sky130_fd_sc_hd__mux2_1
X_14563_ _18390_/Q _14589_/A2 _14589_/B1 input18/X vssd1 vssd1 vccd1 vccd1 _14564_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_260_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11775_ _15039_/B _11774_/X _11726_/B vssd1 vssd1 vccd1 vccd1 _11775_/X sky130_fd_sc_hd__a21o_1
XANTENNA_398 _09457_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _17700_/A0 _18915_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _18915_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _17937_/Q _13742_/A2 _13513_/X _14177_/A vssd1 vssd1 vccd1 vccd1 _17937_/D
+ sky130_fd_sc_hd__o211a_1
X_10726_ _19089_/Q _18993_/Q _10726_/S vssd1 vssd1 vccd1 vccd1 _10726_/X sky130_fd_sc_hd__mux2_1
X_14494_ _17696_/A0 _18344_/Q _14517_/S vssd1 vssd1 vccd1 vccd1 _18344_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17282_ _17280_/Y _17281_/X _16048_/A vssd1 vssd1 vccd1 vccd1 _19444_/D sky130_fd_sc_hd__a21oi_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19021_ _19213_/CLK _19021_/D vssd1 vssd1 vccd1 vccd1 _19021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13445_ _17935_/Q _13742_/A2 _13444_/X _14177_/A vssd1 vssd1 vccd1 vccd1 _17935_/D
+ sky130_fd_sc_hd__o211a_1
X_16233_ _16597_/A0 _18848_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _18848_/D sky130_fd_sc_hd__mux2_1
XFILLER_277_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10657_ _10662_/A1 _19218_/Q _19186_/Q _10656_/S _08899_/A vssd1 vssd1 vccd1 vccd1
+ _10657_/X sky130_fd_sc_hd__a221o_1
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13376_ _19374_/Q _13375_/X _13925_/S vssd1 vssd1 vccd1 vccd1 _13376_/X sky130_fd_sc_hd__mux2_2
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16164_ _16594_/A0 _18781_/Q _16189_/S vssd1 vssd1 vccd1 vccd1 _18781_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10588_ _10586_/X _10587_/X _10663_/S vssd1 vssd1 vccd1 vccd1 _10588_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15115_ _15108_/X _15109_/X _15114_/Y vssd1 vssd1 vccd1 vccd1 _15116_/A sky130_fd_sc_hd__a21oi_2
X_12327_ _17810_/Q _17809_/Q _17808_/Q _17811_/Q vssd1 vssd1 vccd1 vccd1 _12330_/C
+ sky130_fd_sc_hd__or4b_1
X_16095_ _18750_/Q _16095_/B vssd1 vssd1 vccd1 vccd1 _16095_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15046_ _18530_/Q _14666_/X _15045_/X vssd1 vssd1 vccd1 vccd1 _18531_/D sky130_fd_sc_hd__a21oi_1
X_12258_ _17885_/Q _12256_/B _12257_/Y vssd1 vssd1 vccd1 vccd1 _17885_/D sky130_fd_sc_hd__o21a_1
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11209_ _08950_/A _11195_/Y _11208_/X _09523_/A vssd1 vssd1 vccd1 vccd1 _11209_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_269_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189_ _17860_/Q _12192_/C _16768_/A vssd1 vssd1 vccd1 vccd1 _12189_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18805_ _19055_/CLK _18805_/D vssd1 vssd1 vccd1 vccd1 _18805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16997_ _19335_/Q _17043_/B vssd1 vssd1 vccd1 vccd1 _16997_/X sky130_fd_sc_hd__or2_1
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18736_ _18738_/CLK _18736_/D vssd1 vssd1 vccd1 vccd1 _18736_/Q sky130_fd_sc_hd__dfxtp_4
X_15948_ _18691_/Q _15948_/A2 _15948_/B1 _15947_/X _15948_/C1 vssd1 vssd1 vccd1 vccd1
+ _15948_/X sky130_fd_sc_hd__a221o_1
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18667_ _18715_/CLK _18667_/D vssd1 vssd1 vccd1 vccd1 _18667_/Q sky130_fd_sc_hd__dfxtp_1
X_15879_ _18668_/Q _15906_/A2 _15908_/C _15878_/Y _15906_/B1 vssd1 vssd1 vccd1 vccd1
+ _15879_/X sky130_fd_sc_hd__a221o_1
XFILLER_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17618_ _19550_/Q _17624_/A2 _17617_/X _17368_/A vssd1 vssd1 vccd1 vccd1 _19550_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18598_ _19619_/CLK _18598_/D vssd1 vssd1 vccd1 vccd1 _18598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17549_ _17821_/Q _17543_/B1 _17531_/B _13958_/A vssd1 vssd1 vccd1 vccd1 _17550_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_149_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19219_ _19219_/CLK _19219_/D vssd1 vssd1 vccd1 vccd1 _19219_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_93_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18775_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19620_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09805_ _11616_/S _09804_/X _09803_/X _11622_/A1 vssd1 vssd1 vccd1 vccd1 _09805_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09736_ _12999_/S _09736_/B vssd1 vssd1 vccd1 vccd1 _12985_/A sky130_fd_sc_hd__nand2_4
XFILLER_262_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ _18240_/Q _18815_/Q _09671_/S vssd1 vssd1 vccd1 vccd1 _09667_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09598_ _18631_/Q _10717_/S vssd1 vssd1 vccd1 vccd1 _09598_/X sky130_fd_sc_hd__or2_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11560_ _11566_/A1 _19585_/Q _11581_/S _19617_/Q vssd1 vssd1 vccd1 vccd1 _11560_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_126_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10511_ _18868_/Q _18900_/Q _10511_/S vssd1 vssd1 vccd1 vccd1 _10511_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11491_ _18544_/Q _18419_/Q _18028_/Q _17996_/Q _10424_/S _11510_/S1 vssd1 vssd1
+ vccd1 vccd1 _11491_/X sky130_fd_sc_hd__mux4_2
XFILLER_137_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13230_ _12836_/Y _13230_/A1 _13230_/S vssd1 vssd1 vccd1 vccd1 _13230_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10442_ _19644_/Q _18933_/Q _10667_/S vssd1 vssd1 vccd1 vccd1 _10442_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _13201_/B _13161_/B vssd1 vssd1 vccd1 vccd1 _13162_/B sky130_fd_sc_hd__or2_1
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10373_ _10371_/X _10372_/X _10373_/S vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12112_ _17830_/Q _17831_/Q _12112_/C vssd1 vssd1 vccd1 vccd1 _12114_/B sky130_fd_sc_hd__and3_1
XFILLER_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13092_ _13088_/X _13091_/X _13136_/S vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__mux2_2
XFILLER_2_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16920_ _16968_/A _16920_/B vssd1 vssd1 vccd1 vccd1 _19314_/D sky130_fd_sc_hd__and2_1
X_12043_ _16392_/B _12051_/B vssd1 vssd1 vccd1 vccd1 _12043_/X sky130_fd_sc_hd__or2_1
Xfanout1701 _11480_/C1 vssd1 vssd1 vccd1 vccd1 _11397_/A1 sky130_fd_sc_hd__buf_8
Xfanout1712 _08837_/Y vssd1 vssd1 vccd1 vccd1 _09043_/A sky130_fd_sc_hd__buf_6
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1723 _18731_/Q vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1734 _18339_/Q vssd1 vssd1 vccd1 vccd1 _09990_/S sky130_fd_sc_hd__buf_12
XFILLER_172_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16851_ _19297_/Q _16967_/S _16850_/Y _16968_/A vssd1 vssd1 vccd1 vccd1 _19297_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1745 _18202_/Q vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__buf_4
XFILLER_238_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1756 _10689_/S vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__buf_6
XFILLER_93_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1767 _17910_/Q vssd1 vssd1 vccd1 vccd1 _15129_/B2 sky130_fd_sc_hd__clkbuf_16
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1778 _10589_/S vssd1 vssd1 vccd1 vccd1 _11601_/A sky130_fd_sc_hd__buf_6
XFILLER_19_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout780 _16591_/Y vssd1 vssd1 vccd1 vccd1 _16623_/S sky130_fd_sc_hd__buf_8
Xfanout791 _16521_/S vssd1 vssd1 vccd1 vccd1 _16523_/S sky130_fd_sc_hd__buf_12
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15802_ _18594_/Q _16592_/A0 _15817_/S vssd1 vssd1 vccd1 vccd1 _18594_/D sky130_fd_sc_hd__mux2_1
X_19570_ _19602_/CLK _19570_/D vssd1 vssd1 vccd1 vccd1 _19570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1789 _17904_/Q vssd1 vssd1 vccd1 vccd1 _10513_/S sky130_fd_sc_hd__buf_12
X_16782_ _19281_/Q _16783_/C _19282_/Q vssd1 vssd1 vccd1 vccd1 _16784_/B sky130_fd_sc_hd__a21oi_1
X_13994_ _17962_/Q _14032_/B vssd1 vssd1 vccd1 vccd1 _13994_/X sky130_fd_sc_hd__or2_1
XFILLER_253_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18521_ _19286_/CLK _18521_/D vssd1 vssd1 vccd1 vccd1 _18521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _15623_/A _15728_/Y _15732_/Y vssd1 vssd1 vccd1 vccd1 _15733_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _13135_/S _12945_/B vssd1 vssd1 vccd1 vccd1 _12945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18452_ _19631_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _15704_/C _15664_/B vssd1 vssd1 vccd1 vccd1 _15664_/Y sky130_fd_sc_hd__nor2_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12876_ _12674_/X _12695_/X _12943_/S vssd1 vssd1 vccd1 vccd1 _12877_/A sky130_fd_sc_hd__mux2_1
XANTENNA_140 _11836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _11868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_162 _12461_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17403_ _18103_/Q _17437_/A2 _17401_/X _17402_/X vssd1 vssd1 vccd1 vccd1 _17403_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_173 _13998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _16607_/A0 _18422_/Q _14622_/S vssd1 vssd1 vccd1 vccd1 _18422_/D sky130_fd_sc_hd__mux2_1
XANTENNA_184 _13612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11827_ _11899_/A _11827_/B _11827_/C vssd1 vssd1 vccd1 vccd1 _11827_/X sky130_fd_sc_hd__and3_4
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _19399_/CLK _18383_/D vssd1 vssd1 vccd1 vccd1 _18383_/Q sky130_fd_sc_hd__dfxtp_4
X_15595_ _13673_/Y _15110_/X _10750_/Y _15111_/A vssd1 vssd1 vccd1 vccd1 _15595_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_14_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _14030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17334_ _17342_/A _17334_/B vssd1 vssd1 vccd1 vccd1 _19464_/D sky130_fd_sc_hd__and2_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14546_ _14592_/A _14546_/B vssd1 vssd1 vccd1 vccd1 _18381_/D sky130_fd_sc_hd__or2_1
XFILLER_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11758_ _18576_/Q _11759_/A2 _11844_/A _13402_/B vssd1 vssd1 vccd1 vccd1 _11758_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10709_ _09463_/S _10708_/X _09106_/B vssd1 vssd1 vccd1 vccd1 _10709_/X sky130_fd_sc_hd__o21a_1
XFILLER_147_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17265_ _19439_/Q _17310_/B vssd1 vssd1 vccd1 vccd1 _17265_/Y sky130_fd_sc_hd__nand2_1
X_14477_ _18329_/Q _17681_/A0 _14477_/S vssd1 vssd1 vccd1 vccd1 _18329_/D sky130_fd_sc_hd__mux2_1
X_11689_ _11689_/A _14528_/B vssd1 vssd1 vccd1 vccd1 _14525_/A sky130_fd_sc_hd__nand2_8
XFILLER_128_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19004_ _19587_/CLK _19004_/D vssd1 vssd1 vccd1 vccd1 _19004_/Q sky130_fd_sc_hd__dfxtp_1
X_16216_ _17713_/A0 _18832_/Q _16226_/S vssd1 vssd1 vccd1 vccd1 _18832_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13428_ _19537_/Q _13921_/S vssd1 vssd1 vccd1 vccd1 _13428_/X sky130_fd_sc_hd__or2_1
XFILLER_128_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17196_ _17199_/A _17196_/B vssd1 vssd1 vccd1 vccd1 _17517_/A sky130_fd_sc_hd__nand2_1
X_16147_ _18775_/Q _16147_/A2 _16146_/X vssd1 vssd1 vccd1 vccd1 _16154_/B sky130_fd_sc_hd__a21o_1
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13359_ _12835_/A _13353_/X _13356_/X _13602_/B2 _13358_/X vssd1 vssd1 vccd1 vccd1
+ _13359_/X sky130_fd_sc_hd__o221a_1
XFILLER_154_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16078_ _16143_/C _16093_/B _16078_/C vssd1 vssd1 vccd1 vccd1 _16078_/X sky130_fd_sc_hd__or3_4
XFILLER_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15029_ _18518_/Q input195/X _15038_/S vssd1 vssd1 vccd1 vccd1 _18518_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_140_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18272_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_284_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 coreIndex[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_8
XFILLER_49_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09521_ _09978_/A1 _09510_/X _09520_/X _11516_/B1 vssd1 vssd1 vccd1 vccd1 _09521_/X
+ sky130_fd_sc_hd__o211a_1
X_18719_ _18772_/CLK _18719_/D vssd1 vssd1 vccd1 vccd1 _18719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09452_ _18446_/Q _18347_/Q _09464_/S vssd1 vssd1 vccd1 vccd1 _09452_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09383_ _10747_/A1 _09382_/X _09377_/X _11515_/B1 vssd1 vssd1 vccd1 vccd1 _09383_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_212_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput350 _11878_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[24] sky130_fd_sc_hd__buf_4
XFILLER_161_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput361 _11797_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[5] sky130_fd_sc_hd__buf_4
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput372 _11723_/X vssd1 vssd1 vccd1 vccd1 csb0[0] sky130_fd_sc_hd__buf_4
Xoutput383 _11936_/X vssd1 vssd1 vccd1 vccd1 din0[16] sky130_fd_sc_hd__buf_4
XFILLER_266_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1008 _16459_/X vssd1 vssd1 vccd1 vccd1 _16485_/S sky130_fd_sc_hd__buf_12
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput394 _11946_/X vssd1 vssd1 vccd1 vccd1 din0[26] sky130_fd_sc_hd__buf_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1019 _14973_/A1 vssd1 vssd1 vccd1 vccd1 _15003_/A1 sky130_fd_sc_hd__buf_4
XFILLER_102_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09719_ _11190_/A1 _19558_/Q _09720_/S _19590_/Q _09723_/S vssd1 vssd1 vccd1 vccd1
+ _09719_/X sky130_fd_sc_hd__o221a_1
XFILLER_274_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10991_ _19085_/Q _11386_/S _10990_/X _11464_/C1 vssd1 vssd1 vccd1 vccd1 _10991_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _09401_/C _12733_/S _12729_/X vssd1 vssd1 vccd1 vccd1 _12730_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_231_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12656_/A _12659_/Y _12660_/X vssd1 vssd1 vccd1 vccd1 _12661_/X sky130_fd_sc_hd__a21o_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11618_/A1 _19585_/Q _11609_/S _19617_/Q _11616_/S vssd1 vssd1 vccd1 vccd1
+ _11612_/X sky130_fd_sc_hd__o221a_1
X_14400_ _17707_/A0 _18251_/Q _14402_/S vssd1 vssd1 vccd1 vccd1 _18251_/D sky130_fd_sc_hd__mux2_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _15380_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15380_/X sky130_fd_sc_hd__and2_1
X_12592_ _13916_/A _11824_/A _12591_/X vssd1 vssd1 vccd1 vccd1 _12761_/C sky130_fd_sc_hd__o21a_1
XFILLER_129_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11543_ _13727_/A _11642_/B _10603_/A vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__a21o_2
X_14331_ _18188_/Q _17715_/A0 _14339_/S vssd1 vssd1 vccd1 vccd1 _18188_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17050_ _17381_/C _17591_/D vssd1 vssd1 vccd1 vccd1 _17050_/X sky130_fd_sc_hd__or2_4
X_14262_ _18129_/Q _14266_/B vssd1 vssd1 vccd1 vccd1 _14262_/X sky130_fd_sc_hd__or2_1
X_11474_ _09457_/A _11471_/X _11473_/X vssd1 vssd1 vccd1 vccd1 _11474_/Y sky130_fd_sc_hd__a21oi_2
X_16001_ _18716_/Q _16005_/A2 _16000_/X _14205_/A vssd1 vssd1 vccd1 vccd1 _18716_/D
+ sky130_fd_sc_hd__o211a_1
X_13213_ _19369_/Q _13951_/A2 _13211_/X _13212_/X _13951_/C1 vssd1 vssd1 vccd1 vccd1
+ _13213_/X sky130_fd_sc_hd__o221a_4
X_10425_ _10427_/C1 _10424_/X _10423_/X _11503_/S1 vssd1 vssd1 vccd1 vccd1 _10425_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14193_ _16964_/A _14193_/B vssd1 vssd1 vccd1 vccd1 _18094_/D sky130_fd_sc_hd__and2_1
XFILLER_125_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13144_ _12448_/D _13128_/X _13143_/Y _13124_/X vssd1 vssd1 vccd1 vccd1 _13144_/X
+ sky130_fd_sc_hd__a31o_1
X_10356_ _10200_/S _10348_/X _10347_/X _10356_/C1 vssd1 vssd1 vccd1 vccd1 _10356_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_11__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_78_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13075_ _13945_/B2 _13059_/X _13074_/X vssd1 vssd1 vccd1 vccd1 _13986_/B sky130_fd_sc_hd__a21oi_4
X_17952_ _18627_/CLK _17952_/D vssd1 vssd1 vccd1 vccd1 _17952_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10287_ _19063_/Q _19031_/Q _10299_/S vssd1 vssd1 vccd1 vccd1 _10287_/X sky130_fd_sc_hd__mux2_1
XFILLER_250_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1520 _10426_/S vssd1 vssd1 vccd1 vccd1 _11513_/B2 sky130_fd_sc_hd__buf_6
XFILLER_239_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16903_ _19310_/Q _17587_/A _16971_/S vssd1 vssd1 vccd1 vccd1 _16904_/B sky130_fd_sc_hd__mux2_1
X_12026_ _17888_/Q _12052_/A2 _12025_/X _13257_/A vssd1 vssd1 vccd1 vccd1 _17790_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1531 _11189_/A vssd1 vssd1 vccd1 vccd1 _10719_/S sky130_fd_sc_hd__buf_4
X_17883_ _19261_/CLK _17883_/D vssd1 vssd1 vccd1 vccd1 _17883_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1542 _11606_/S vssd1 vssd1 vccd1 vccd1 _11355_/A1 sky130_fd_sc_hd__buf_6
XFILLER_266_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1553 _10280_/S vssd1 vssd1 vccd1 vccd1 _09972_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_78_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1564 _11515_/B1 vssd1 vssd1 vccd1 vccd1 _11501_/B1 sky130_fd_sc_hd__buf_8
X_19622_ _19622_/CLK _19622_/D vssd1 vssd1 vccd1 vccd1 _19622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16834_ _17051_/B _17051_/C vssd1 vssd1 vccd1 vccd1 _16975_/B sky130_fd_sc_hd__or2_1
Xfanout1575 fanout1581/X vssd1 vssd1 vccd1 vccd1 _11198_/S sky130_fd_sc_hd__buf_8
Xfanout1586 _10211_/A1 vssd1 vssd1 vccd1 vccd1 _11274_/S1 sky130_fd_sc_hd__buf_6
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1597 _08893_/Y vssd1 vssd1 vccd1 vccd1 _11621_/C1 sky130_fd_sc_hd__clkbuf_16
XFILLER_238_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19553_ _19553_/CLK _19553_/D vssd1 vssd1 vccd1 vccd1 _19553_/Q sky130_fd_sc_hd__dfxtp_1
X_16765_ _19275_/Q _16767_/C _16764_/Y vssd1 vssd1 vccd1 vccd1 _19275_/D sky130_fd_sc_hd__a21oi_1
XFILLER_253_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13977_ _17953_/Q _14034_/B _13976_/Y _14001_/C1 vssd1 vssd1 vccd1 vccd1 _17953_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18504_ _19229_/CLK _18504_/D vssd1 vssd1 vccd1 vccd1 _18504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15716_ _19483_/Q _15715_/Y _15716_/S vssd1 vssd1 vccd1 vccd1 _15716_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19484_ _19484_/CLK _19484_/D vssd1 vssd1 vccd1 vccd1 _19484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _13421_/A _12956_/A _12761_/B _12927_/Y _13185_/A vssd1 vssd1 vccd1 vccd1
+ _12928_/X sky130_fd_sc_hd__a221o_1
X_16696_ _16795_/A _16696_/B _16697_/B vssd1 vssd1 vccd1 vccd1 _19251_/D sky130_fd_sc_hd__nor3_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18435_ _19614_/CLK _18435_/D vssd1 vssd1 vccd1 vccd1 _18435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15647_ _08819_/Y _15751_/A _15731_/B1 _15646_/Y _15717_/B2 vssd1 vssd1 vccd1 vccd1
+ _15647_/X sky130_fd_sc_hd__a221o_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _12851_/X _12858_/X _12859_/S vssd1 vssd1 vccd1 vccd1 _12859_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18366_ _19644_/CLK _18366_/D vssd1 vssd1 vccd1 vccd1 _18366_/Q sky130_fd_sc_hd__dfxtp_1
X_15578_ _15787_/A _15639_/A vssd1 vssd1 vccd1 vccd1 _15638_/B sky130_fd_sc_hd__xnor2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17317_ _19456_/Q _17117_/B _17377_/S vssd1 vssd1 vccd1 vccd1 _17318_/B sky130_fd_sc_hd__mux2_1
X_14529_ _18373_/Q _14575_/A2 _14575_/B1 input10/X vssd1 vssd1 vccd1 vccd1 _14530_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18297_ _19450_/CLK _18297_/D vssd1 vssd1 vccd1 vccd1 _18297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17248_ _14224_/A _17166_/A _17438_/A _17310_/B vssd1 vssd1 vccd1 vccd1 _17248_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_179_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17179_ _19411_/Q fanout533/X _17488_/A _17120_/B vssd1 vssd1 vccd1 vccd1 _17180_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_190_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ _11508_/B1 _14306_/C _16459_/A _10217_/B _08950_/Y vssd1 vssd1 vccd1 vccd1
+ _08956_/C sky130_fd_sc_hd__o221a_1
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08883_ _08883_/A vssd1 vssd1 vccd1 vccd1 _08883_/Y sky130_fd_sc_hd__inv_6
XFILLER_229_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09504_ _09502_/X _09503_/X _09972_/S vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09435_ _11055_/B2 _09432_/X _09437_/B _11210_/A1 vssd1 vssd1 vccd1 vccd1 _15238_/A
+ sky130_fd_sc_hd__a2bb2o_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09366_ _17916_/Q _09140_/S _09367_/B vssd1 vssd1 vccd1 vccd1 _09401_/B sky130_fd_sc_hd__o21ai_4
XFILLER_240_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09297_ _08896_/A _09296_/X _09289_/X _11501_/B1 vssd1 vssd1 vccd1 vccd1 _09297_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_40 _11812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_51 _12613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_62 _13917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_73 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_84 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_95 _11845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10210_ _11046_/S1 _10200_/X _10209_/X _11438_/B1 vssd1 vssd1 vccd1 vccd1 _10210_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ _11190_/A1 _18955_/Q _18220_/Q _09883_/B vssd1 vssd1 vccd1 vccd1 _11190_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10141_ _18624_/Q _18195_/Q _10141_/S vssd1 vssd1 vccd1 vccd1 _10141_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10072_ _11739_/A _11739_/B _13044_/S vssd1 vssd1 vccd1 vccd1 _11743_/A sky130_fd_sc_hd__a21oi_4
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13900_ _18130_/Q _18129_/Q _13900_/C vssd1 vssd1 vccd1 vccd1 _13934_/B sky130_fd_sc_hd__and3_2
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14880_ _18489_/Q _15001_/A2 _14879_/Y _16795_/A vssd1 vssd1 vccd1 vccd1 _18489_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_208_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13831_ _14028_/B vssd1 vssd1 vccd1 vccd1 _13831_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16550_ _10532_/B _19155_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _19155_/D sky130_fd_sc_hd__mux2_1
X_13762_ _10604_/Y _13727_/B _12650_/X vssd1 vssd1 vccd1 vccd1 _13763_/B sky130_fd_sc_hd__a21oi_2
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10974_ _11355_/A1 _10973_/X _11623_/A1 vssd1 vssd1 vccd1 vccd1 _10974_/X sky130_fd_sc_hd__a21o_1
XFILLER_204_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _17906_/Q _15452_/A _15484_/A vssd1 vssd1 vccd1 vccd1 _15506_/A sky130_fd_sc_hd__o21ai_2
XFILLER_71_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12713_ _12712_/X _12711_/X _12813_/S vssd1 vssd1 vccd1 vccd1 _12713_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16481_ _16547_/A0 _19088_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _19088_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13693_ _13930_/A1 _13679_/Y _13930_/B1 vssd1 vssd1 vccd1 vccd1 _13693_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18220_ _19147_/CLK _18220_/D vssd1 vssd1 vccd1 vccd1 _18220_/Q sky130_fd_sc_hd__dfxtp_1
X_15432_ _15432_/A _15432_/B vssd1 vssd1 vccd1 vccd1 _15456_/D sky130_fd_sc_hd__xnor2_2
X_12644_ _12639_/Y _12643_/Y _13697_/A vssd1 vssd1 vccd1 vccd1 _12644_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_231_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18151_ _19047_/CLK _18151_/D vssd1 vssd1 vccd1 vccd1 _18151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12575_ _12575_/A _12584_/B vssd1 vssd1 vccd1 vccd1 _12575_/Y sky130_fd_sc_hd__nor2_8
X_15363_ _15310_/A _15308_/B _15362_/X _15335_/X _15306_/Y vssd1 vssd1 vccd1 vccd1
+ _15364_/B sky130_fd_sc_hd__a311o_2
X_17102_ _17193_/B _17108_/A2 _17101_/X _17366_/A vssd1 vssd1 vccd1 vccd1 _19384_/D
+ sky130_fd_sc_hd__o211a_1
X_14314_ _18171_/Q _15808_/A1 _14335_/S vssd1 vssd1 vccd1 vccd1 _18171_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18082_ _19304_/CLK _18082_/D vssd1 vssd1 vccd1 vccd1 _18082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11526_ _11681_/A _11681_/B _13316_/A vssd1 vssd1 vccd1 vccd1 _11680_/B sky130_fd_sc_hd__o21bai_4
XFILLER_129_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15294_ _12788_/B _15293_/X _15307_/B vssd1 vssd1 vccd1 vccd1 _15294_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17033_ _19353_/Q _17041_/B vssd1 vssd1 vccd1 vccd1 _17033_/X sky130_fd_sc_hd__or2_1
X_11457_ _11465_/A1 _18216_/Q _11462_/S _18951_/Q _11464_/C1 vssd1 vssd1 vccd1 vccd1
+ _11457_/X sky130_fd_sc_hd__o221a_1
XFILLER_172_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14245_ _18294_/Q _14267_/A2 _14244_/X _14442_/B vssd1 vssd1 vccd1 vccd1 _18120_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10408_ _10406_/X _10407_/X _10408_/S vssd1 vssd1 vccd1 vccd1 _10409_/B sky130_fd_sc_hd__mux2_1
XFILLER_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14176_ _18699_/Q _18086_/Q _14186_/S vssd1 vssd1 vccd1 vccd1 _14177_/B sky130_fd_sc_hd__mux2_1
XFILLER_171_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11388_ _11389_/A1 _19567_/Q _11384_/B _19599_/Q _11464_/C1 vssd1 vssd1 vccd1 vccd1
+ _11388_/X sky130_fd_sc_hd__o221a_1
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _10336_/X _10338_/X _10332_/X vssd1 vssd1 vccd1 vccd1 _10339_/Y sky130_fd_sc_hd__a21oi_4
X_13127_ _13127_/A _13127_/B vssd1 vssd1 vccd1 vccd1 _14143_/A sky130_fd_sc_hd__xnor2_2
X_18984_ _19565_/CLK _18984_/D vssd1 vssd1 vccd1 vccd1 _18984_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _18660_/CLK _17935_/D vssd1 vssd1 vccd1 vccd1 _17935_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _15214_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _13058_/X sky130_fd_sc_hd__or2_1
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12009_ _17776_/Q _17677_/A0 _12021_/S vssd1 vssd1 vccd1 vccd1 _17776_/D sky130_fd_sc_hd__mux2_1
Xfanout1350 _09919_/C1 vssd1 vssd1 vccd1 vccd1 _10250_/S sky130_fd_sc_hd__buf_8
XFILLER_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1361 _11167_/B vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__buf_6
XFILLER_39_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17866_ _19327_/CLK _17866_/D vssd1 vssd1 vccd1 vccd1 _17866_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1372 _10613_/S vssd1 vssd1 vccd1 vccd1 _10619_/S sky130_fd_sc_hd__buf_6
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1383 fanout1386/X vssd1 vssd1 vccd1 vccd1 _11249_/S sky130_fd_sc_hd__buf_6
Xfanout1394 _10320_/S vssd1 vssd1 vccd1 vccd1 _09688_/S sky130_fd_sc_hd__buf_4
XFILLER_281_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16817_ _08821_/Y _16816_/C _16964_/A vssd1 vssd1 vccd1 vccd1 _16817_/Y sky130_fd_sc_hd__o21ai_1
X_19605_ _19632_/CLK _19605_/D vssd1 vssd1 vccd1 vccd1 _19605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17797_ _18201_/CLK _17797_/D vssd1 vssd1 vccd1 vccd1 _17797_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_226_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19536_ _19552_/CLK _19536_/D vssd1 vssd1 vccd1 vccd1 _19536_/Q sky130_fd_sc_hd__dfxtp_1
X_16748_ _19269_/Q _16751_/C _16780_/B1 vssd1 vssd1 vccd1 vccd1 _16748_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_253_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19467_ _19502_/CLK _19467_/D vssd1 vssd1 vccd1 vccd1 _19467_/Q sky130_fd_sc_hd__dfxtp_4
X_16679_ _17724_/A _19246_/Q _19242_/Q _19238_/Q vssd1 vssd1 vccd1 vccd1 _16680_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_146_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ _10346_/S _09218_/X _09219_/X _10356_/C1 vssd1 vssd1 vccd1 vccd1 _09220_/X
+ sky130_fd_sc_hd__a211o_1
X_18418_ _18543_/CLK _18418_/D vssd1 vssd1 vccd1 vccd1 _18418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19398_ _19533_/CLK _19398_/D vssd1 vssd1 vccd1 vccd1 _19398_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ _09034_/B _09150_/X _09326_/A vssd1 vssd1 vccd1 vccd1 _09151_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18349_ _19627_/CLK _18349_/D vssd1 vssd1 vccd1 vccd1 _18349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09082_ _11706_/C _13622_/A vssd1 vssd1 vccd1 vccd1 _15081_/A sky130_fd_sc_hd__nor2_8
XFILLER_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput60 dout0[25] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput71 dout0[35] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_2
Xinput82 dout0[45] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_2
Xinput93 dout0[55] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09984_ _09984_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _12842_/A sky130_fd_sc_hd__xor2_4
XFILLER_131_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08935_ _17821_/Q _17815_/Q _08935_/C vssd1 vssd1 vccd1 vccd1 _08935_/X sky130_fd_sc_hd__or3_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08866_ _17889_/Q _17888_/Q _09062_/B vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__nand3_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09418_ _18633_/Q _18055_/Q _19074_/Q _18978_/Q _09704_/S _11199_/S1 vssd1 vssd1
+ vccd1 vccd1 _09419_/B sky130_fd_sc_hd__mux4_1
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ _18258_/Q _18833_/Q _11249_/S vssd1 vssd1 vccd1 vccd1 _10690_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09349_ _10262_/A1 _18602_/Q _18173_/Q _11481_/C vssd1 vssd1 vccd1 vccd1 _09349_/X
+ sky130_fd_sc_hd__a22o_1
X_12360_ _17895_/Q _12382_/A vssd1 vssd1 vccd1 vccd1 _12360_/X sky130_fd_sc_hd__or2_1
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11311_ _11572_/A1 _19568_/Q _10940_/S _19600_/Q _11311_/C1 vssd1 vssd1 vccd1 vccd1
+ _11311_/X sky130_fd_sc_hd__o221a_1
X_12291_ _14682_/A _12292_/C vssd1 vssd1 vccd1 vccd1 _14679_/B sky130_fd_sc_hd__nor2_1
XFILLER_181_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14030_ _14032_/B _14030_/B vssd1 vssd1 vccd1 vccd1 _14030_/Y sky130_fd_sc_hd__nand2_1
X_11242_ _11251_/S _19178_/Q _11247_/S vssd1 vssd1 vccd1 vccd1 _11242_/X sky130_fd_sc_hd__and3_1
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11173_ _11171_/X _11172_/X _11173_/S vssd1 vssd1 vccd1 vccd1 _11173_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10124_ _18562_/Q _18437_/Q _10206_/S vssd1 vssd1 vccd1 vccd1 _10124_/X sky130_fd_sc_hd__mux2_1
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15981_ _18706_/Q _16019_/A2 _15980_/X _16964_/A vssd1 vssd1 vccd1 vccd1 _18706_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _17720_/A0 _19646_/Q _17722_/S vssd1 vssd1 vccd1 vccd1 _19646_/D sky130_fd_sc_hd__mux2_1
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10055_ _11618_/A1 _18204_/Q _11617_/S _18939_/Q _10745_/S vssd1 vssd1 vccd1 vccd1
+ _10055_/X sky130_fd_sc_hd__o221a_1
X_14932_ _15003_/A1 _13723_/X _15003_/B1 _18650_/Q _15003_/C1 vssd1 vssd1 vccd1 vccd1
+ _14932_/X sky130_fd_sc_hd__a221o_1
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17651_ _17684_/A0 _19579_/Q _17657_/S vssd1 vssd1 vccd1 vccd1 _19579_/D sky130_fd_sc_hd__mux2_1
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ _14861_/X _14862_/X _14714_/B vssd1 vssd1 vccd1 vccd1 _14863_/X sky130_fd_sc_hd__a21o_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ _16602_/A0 _19205_/Q _16622_/S vssd1 vssd1 vccd1 vccd1 _19205_/D sky130_fd_sc_hd__mux2_1
X_13814_ _10380_/Y _13912_/B1 _13912_/A2 _11550_/B _14153_/A vssd1 vssd1 vccd1 vccd1
+ _13814_/X sky130_fd_sc_hd__a221o_1
XFILLER_217_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17582_ _19533_/Q _17558_/B _17603_/B1 _17581_/X vssd1 vssd1 vccd1 vccd1 _19533_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_235_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14794_ input44/X input79/X _14844_/S vssd1 vssd1 vccd1 vccd1 _14795_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19321_ _19321_/CLK _19321_/D vssd1 vssd1 vccd1 vccd1 _19321_/Q sky130_fd_sc_hd__dfxtp_1
X_16533_ _09437_/B _19138_/Q _16554_/S vssd1 vssd1 vccd1 vccd1 _19138_/D sky130_fd_sc_hd__mux2_1
X_13745_ _19257_/Q _13943_/A2 _13943_/B1 _19289_/Q vssd1 vssd1 vccd1 vccd1 _13745_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10957_ _18645_/Q _18067_/Q _19086_/Q _18990_/Q _11613_/S _11338_/S1 vssd1 vssd1
+ vccd1 vccd1 _10958_/B sky130_fd_sc_hd__mux4_1
XFILLER_32_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19252_ _19261_/CLK _19252_/D vssd1 vssd1 vccd1 vccd1 _19252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16464_ _17663_/A0 _19071_/Q _16485_/S vssd1 vssd1 vccd1 vccd1 _19071_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13676_ _13938_/A _13676_/B vssd1 vssd1 vccd1 vccd1 _13676_/Y sky130_fd_sc_hd__nand2_1
X_10888_ _11596_/A1 _19215_/Q _19183_/Q _10815_/B vssd1 vssd1 vccd1 vccd1 _10888_/X
+ sky130_fd_sc_hd__a22o_1
X_18203_ _19650_/CLK _18203_/D vssd1 vssd1 vccd1 vccd1 _18203_/Q sky130_fd_sc_hd__dfxtp_1
X_15415_ _15789_/A1 _15410_/Y _15437_/B1 vssd1 vssd1 vccd1 vccd1 _15416_/C sky130_fd_sc_hd__a21oi_2
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19183_ _19607_/CLK _19183_/D vssd1 vssd1 vccd1 vccd1 _19183_/Q sky130_fd_sc_hd__dfxtp_1
X_12627_ _12624_/A _12624_/B _12626_/X vssd1 vssd1 vccd1 vccd1 _13465_/B sky130_fd_sc_hd__a21o_2
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16395_ _16593_/A0 _19004_/Q _16424_/S vssd1 vssd1 vccd1 vccd1 _19004_/D sky130_fd_sc_hd__mux2_1
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18134_ _19619_/CLK _18134_/D vssd1 vssd1 vccd1 vccd1 _18134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15346_ _15319_/Y _15324_/B _15321_/B vssd1 vssd1 vccd1 vccd1 _15347_/B sky130_fd_sc_hd__o21ai_2
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _13167_/A _12561_/B vssd1 vssd1 vccd1 vccd1 _12558_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11509_ _11509_/A _11509_/B vssd1 vssd1 vccd1 vccd1 _11509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18065_ _19134_/CLK _18065_/D vssd1 vssd1 vccd1 vccd1 _18065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15277_ _15275_/Y _15277_/B vssd1 vssd1 vccd1 vccd1 _15280_/A sky130_fd_sc_hd__nand2b_1
X_12489_ _12488_/A _14682_/A _12488_/Y vssd1 vssd1 vccd1 vccd1 _12572_/C sky130_fd_sc_hd__o21ai_2
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17016_ _17169_/B _17032_/A2 _17015_/X _17360_/A vssd1 vssd1 vccd1 vccd1 _19344_/D
+ sky130_fd_sc_hd__o211a_1
X_14228_ _18112_/Q _14266_/B vssd1 vssd1 vccd1 vccd1 _14228_/X sky130_fd_sc_hd__or2_1
XFILLER_171_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ _12263_/A _15328_/C _12461_/A vssd1 vssd1 vccd1 vccd1 _14159_/Y sky130_fd_sc_hd__o21ai_2
Xfanout609 _12571_/X vssd1 vssd1 vccd1 vccd1 _13247_/C1 sky130_fd_sc_hd__buf_6
XFILLER_217_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18967_ _19159_/CLK _18967_/D vssd1 vssd1 vccd1 vccd1 _18967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17918_ _19595_/CLK _17918_/D vssd1 vssd1 vccd1 vccd1 _17918_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_47_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19625_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_239_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18898_ _19641_/CLK _18898_/D vssd1 vssd1 vccd1 vccd1 _18898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_255_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1180 _15526_/B vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__buf_4
XFILLER_254_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1191 _16004_/B1 vssd1 vssd1 vccd1 vccd1 _16147_/A2 sky130_fd_sc_hd__buf_4
X_17849_ _19324_/CLK _17849_/D vssd1 vssd1 vccd1 vccd1 _17849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19519_ _19519_/CLK _19519_/D vssd1 vssd1 vccd1 vccd1 _19519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09203_ _09708_/A _09203_/B vssd1 vssd1 vccd1 vccd1 _09203_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09134_ _18950_/Q _18215_/Q _11455_/S vssd1 vssd1 vccd1 vccd1 _09134_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09065_ _17900_/Q _12665_/B vssd1 vssd1 vccd1 vccd1 _11647_/A sky130_fd_sc_hd__or2_4
XFILLER_108_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ _09965_/X _09966_/X _09967_/S vssd1 vssd1 vccd1 vccd1 _09967_/X sky130_fd_sc_hd__mux2_1
XFILLER_246_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08918_ _12089_/A _17800_/Q vssd1 vssd1 vccd1 vccd1 _14488_/C sky130_fd_sc_hd__and2_2
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09898_/A _12602_/B vssd1 vssd1 vccd1 vccd1 _11731_/B sky130_fd_sc_hd__nand2_2
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08849_ _10036_/S vssd1 vssd1 vccd1 vccd1 _08849_/Y sky130_fd_sc_hd__inv_2
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_503 _10027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_514 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _11860_/A _11864_/B vssd1 vssd1 vccd1 vccd1 _11896_/A sky130_fd_sc_hd__or2_2
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_525 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_536 input225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _18615_/Q _18186_/Q _11598_/S vssd1 vssd1 vccd1 vccd1 _10811_/X sky130_fd_sc_hd__mux2_1
XANTENNA_547 _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11791_ _11820_/A wire989/X vssd1 vssd1 vccd1 vccd1 _11791_/Y sky130_fd_sc_hd__nand2_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13530_ _13791_/A _13528_/X _13529_/Y _13545_/B _13622_/A vssd1 vssd1 vccd1 vccd1
+ _13530_/X sky130_fd_sc_hd__a32o_1
X_10742_ _10742_/A1 _10734_/X _10735_/X vssd1 vssd1 vccd1 vccd1 _10742_/X sky130_fd_sc_hd__o21a_1
XFILLER_213_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10673_ _11365_/B2 _16615_/A0 _10672_/X _11133_/B2 vssd1 vssd1 vccd1 vccd1 _13679_/A
+ sky130_fd_sc_hd__o2bb2a_4
X_13461_ _12586_/X _13446_/Y _13563_/B1 vssd1 vssd1 vccd1 vccd1 _13462_/C sky130_fd_sc_hd__a21o_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ _15200_/A _15200_/B vssd1 vssd1 vccd1 vccd1 _15207_/B sky130_fd_sc_hd__nor2_1
X_12412_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12412_/Y sky130_fd_sc_hd__nand2_1
X_16180_ _16610_/A0 _18797_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _18797_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13392_ _11369_/A _13316_/B _14156_/A0 vssd1 vssd1 vccd1 vccd1 _13392_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15131_ _15259_/B _12869_/Y _15285_/A3 _15130_/X vssd1 vssd1 vccd1 vccd1 _15131_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_182_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12343_ _12349_/A _12343_/B vssd1 vssd1 vccd1 vccd1 _12343_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12274_ _18776_/Q _18775_/Q vssd1 vssd1 vccd1 vccd1 _16095_/B sky130_fd_sc_hd__or2_4
X_15062_ _18546_/Q _16540_/A0 _15079_/S vssd1 vssd1 vccd1 vccd1 _18546_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14013_ _17971_/Q _14020_/B _14012_/Y _14037_/C1 vssd1 vssd1 vccd1 vccd1 _17971_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11225_ _19082_/Q _11226_/S _11224_/X _11569_/S1 vssd1 vssd1 vccd1 vccd1 _11225_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18821_ _19126_/CLK _18821_/D vssd1 vssd1 vccd1 vccd1 _18821_/Q sky130_fd_sc_hd__dfxtp_1
X_11156_ _11157_/A1 _19570_/Q _11154_/S _19602_/Q _11156_/C1 vssd1 vssd1 vccd1 vccd1
+ _11156_/X sky130_fd_sc_hd__o221a_1
XFILLER_110_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10107_ _10334_/A1 _19584_/Q _10090_/S _19616_/Q vssd1 vssd1 vccd1 vccd1 _10107_/X
+ sky130_fd_sc_hd__o22a_1
X_18752_ _18776_/CLK _18752_/D vssd1 vssd1 vccd1 vccd1 _18752_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15964_ _18697_/Q _15970_/A2 _15976_/B1 _18746_/Q _15976_/C1 vssd1 vssd1 vccd1 vccd1
+ _15964_/X sky130_fd_sc_hd__a221o_1
X_11087_ _19212_/Q _11482_/A2 _11086_/X _11578_/S vssd1 vssd1 vccd1 vccd1 _11087_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_249_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput250 localMemory_wb_sel_i[3] vssd1 vssd1 vccd1 vccd1 input250/X sky130_fd_sc_hd__clkbuf_2
Xinput261 manufacturerID[7] vssd1 vssd1 vccd1 vccd1 input261/X sky130_fd_sc_hd__clkbuf_4
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17703_ _17703_/A0 _19629_/Q _17722_/S vssd1 vssd1 vccd1 vccd1 _19629_/D sky130_fd_sc_hd__mux2_1
XFILLER_236_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput272 partID[2] vssd1 vssd1 vccd1 vccd1 input272/X sky130_fd_sc_hd__clkbuf_2
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14915_ _15006_/A1 _14914_/X _15006_/B1 vssd1 vssd1 vccd1 vccd1 _14915_/Y sky130_fd_sc_hd__o21ai_2
X_10038_ _18439_/Q _18340_/Q _11613_/S vssd1 vssd1 vccd1 vccd1 _10038_/X sky130_fd_sc_hd__mux2_1
Xinput283 versionID[3] vssd1 vssd1 vccd1 vccd1 input283/X sky130_fd_sc_hd__buf_2
X_18683_ _18683_/CLK _18683_/D vssd1 vssd1 vccd1 vccd1 _18683_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15895_ _18674_/Q _15910_/A2 _15894_/X _15904_/C1 vssd1 vssd1 vccd1 vccd1 _18674_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17634_ _17667_/A0 _19562_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _19562_/D sky130_fd_sc_hd__mux2_1
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ _14696_/A _18270_/Q _14845_/Y _14846_/B1 vssd1 vssd1 vccd1 vccd1 _14846_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17565_ _17589_/B _17565_/B vssd1 vssd1 vccd1 vccd1 _17565_/Y sky130_fd_sc_hd__nand2b_1
X_14777_ _14773_/Y _14776_/X _14879_/B1 vssd1 vssd1 vccd1 vccd1 _14777_/Y sky130_fd_sc_hd__a21oi_4
X_11989_ _17800_/Q _16392_/B _14488_/B vssd1 vssd1 vccd1 vccd1 _14599_/A sky130_fd_sc_hd__or3_4
XFILLER_205_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19304_ _19304_/CLK _19304_/D vssd1 vssd1 vccd1 vccd1 _19304_/Q sky130_fd_sc_hd__dfxtp_1
X_16516_ _16549_/A0 _19122_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _19122_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13728_ _13761_/B _14148_/B _13892_/B1 vssd1 vssd1 vccd1 vccd1 _13728_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_210_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17496_ _18583_/Q _17544_/A _08883_/A vssd1 vssd1 vccd1 vccd1 _17496_/X sky130_fd_sc_hd__o21a_1
XFILLER_220_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_165_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19483_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19235_ _19268_/CLK _19235_/D vssd1 vssd1 vccd1 vccd1 _19235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16447_ _19055_/Q _17712_/A0 _16453_/S vssd1 vssd1 vccd1 vccd1 _19055_/D sky130_fd_sc_hd__mux2_1
XFILLER_220_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13659_ _13649_/Y _13658_/Y _13682_/B2 _13648_/X vssd1 vssd1 vccd1 vccd1 _13659_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19166_ _19621_/CLK _19166_/D vssd1 vssd1 vccd1 vccd1 _19166_/Q sky130_fd_sc_hd__dfxtp_1
X_16378_ _17677_/A0 _18989_/Q _16390_/S vssd1 vssd1 vccd1 vccd1 _18989_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18117_ _18593_/CLK _18117_/D vssd1 vssd1 vccd1 vccd1 _18117_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15329_ _15549_/A _15329_/B vssd1 vssd1 vccd1 vccd1 _15330_/B sky130_fd_sc_hd__nor2_2
X_19097_ _19126_/CLK _19097_/D vssd1 vssd1 vccd1 vccd1 _19097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18048_ _19195_/CLK _18048_/D vssd1 vssd1 vccd1 vccd1 _18048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09821_ _09821_/A _09821_/B _09156_/X vssd1 vssd1 vccd1 vccd1 _09821_/X sky130_fd_sc_hd__or3b_2
XFILLER_63_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09752_ _19006_/Q _11224_/B _09751_/X _09095_/A vssd1 vssd1 vccd1 vccd1 _09752_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_274_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09683_ _09683_/A _09683_/B vssd1 vssd1 vccd1 vccd1 _09683_/X sky130_fd_sc_hd__or2_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09117_ _12468_/B _19206_/Q _19174_/Q _09925_/S _09683_/A vssd1 vssd1 vccd1 vccd1
+ _09117_/X sky130_fd_sc_hd__a221o_1
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ _09048_/A _09331_/A vssd1 vssd1 vccd1 vccd1 _09050_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _11397_/A1 _11007_/X _11008_/X _11009_/X vssd1 vssd1 vccd1 vccd1 _11010_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1905 _14487_/A vssd1 vssd1 vccd1 vccd1 fanout1905/X sky130_fd_sc_hd__buf_8
XFILLER_277_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout940 _14973_/C1 vssd1 vssd1 vccd1 vccd1 _14741_/B sky130_fd_sc_hd__buf_4
XFILLER_77_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout951 _14648_/S vssd1 vssd1 vccd1 vccd1 _14660_/S sky130_fd_sc_hd__buf_12
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout962 _14108_/Y vssd1 vssd1 vccd1 vccd1 _14131_/S sky130_fd_sc_hd__buf_8
XFILLER_265_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout973 _13747_/B2 vssd1 vssd1 vccd1 vccd1 _13682_/B2 sky130_fd_sc_hd__buf_6
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout984 _13808_/C1 vssd1 vssd1 vccd1 vccd1 _13256_/B1 sky130_fd_sc_hd__buf_4
XFILLER_218_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 _10531_/X vssd1 vssd1 vccd1 vccd1 _10532_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_218_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _13100_/A _12961_/B vssd1 vssd1 vccd1 vccd1 _17923_/D sky130_fd_sc_hd__and2_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _14720_/A _14700_/B vssd1 vssd1 vccd1 vccd1 _14700_/Y sky130_fd_sc_hd__nor2_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11912_ _18566_/Q _11663_/A _11706_/B _11737_/X vssd1 vssd1 vccd1 vccd1 _11912_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_246_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _13804_/X _15110_/X _10450_/Y _15111_/A vssd1 vssd1 vccd1 vccd1 _15680_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_300 _18737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ _09897_/Y _14155_/B _13358_/A1 vssd1 vssd1 vccd1 vccd1 _12892_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_311 _18114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_322 _18107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14631_ _17690_/A0 _18438_/Q _14631_/S vssd1 vssd1 vccd1 vccd1 _18438_/D sky130_fd_sc_hd__mux2_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _11952_/A2 _11841_/X _11842_/X vssd1 vssd1 vccd1 vccd1 _11844_/B sky130_fd_sc_hd__a21oi_4
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 _11479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_355 _12461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_366 _08874_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_377 _14889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17350_ _17350_/A _17350_/B vssd1 vssd1 vccd1 vccd1 _19472_/D sky130_fd_sc_hd__and2_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_388 _17003_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14562_ _14586_/A _14562_/B vssd1 vssd1 vccd1 vccd1 _18389_/D sky130_fd_sc_hd__or2_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11774_ _11810_/A _11774_/B _11779_/B vssd1 vssd1 vccd1 vccd1 _11774_/X sky130_fd_sc_hd__and3_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_399 _12609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _17699_/A0 _18914_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _18914_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13513_ _08874_/D _13971_/A2 _13511_/Y _13512_/X _13579_/A vssd1 vssd1 vccd1 vccd1
+ _13513_/X sky130_fd_sc_hd__a221o_4
X_10725_ _10745_/S _10724_/X _10723_/X _11622_/A1 vssd1 vssd1 vccd1 vccd1 _10725_/X
+ sky130_fd_sc_hd__a211o_1
X_17281_ _18121_/Q _17540_/B1 _17493_/A _17289_/B vssd1 vssd1 vccd1 vccd1 _17281_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _17695_/A0 _18343_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _18343_/D sky130_fd_sc_hd__mux2_1
X_19020_ _19621_/CLK _19020_/D vssd1 vssd1 vccd1 vccd1 _19020_/Q sky130_fd_sc_hd__dfxtp_1
X_16232_ _16431_/A1 _18847_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _18847_/D sky130_fd_sc_hd__mux2_1
X_13444_ _09494_/A _12448_/C _13442_/Y _13443_/X _12762_/B vssd1 vssd1 vccd1 vccd1
+ _13444_/X sky130_fd_sc_hd__a221o_4
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10656_ _19058_/Q _19026_/Q _10656_/S vssd1 vssd1 vccd1 vccd1 _10656_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16163_ _17693_/A0 _18780_/Q _16165_/S vssd1 vssd1 vccd1 vccd1 _18780_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13375_ _19470_/Q _12529_/Y _12578_/Y _19342_/Q _13374_/X vssd1 vssd1 vccd1 vccd1
+ _13375_/X sky130_fd_sc_hd__a221o_1
X_10587_ _10662_/A1 _18157_/Q _18803_/Q _10656_/S vssd1 vssd1 vccd1 vccd1 _10587_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15114_ _15108_/X _15369_/A _15109_/X vssd1 vssd1 vccd1 vccd1 _15114_/Y sky130_fd_sc_hd__a21oi_1
X_12326_ _17800_/Q _16392_/B _17798_/Q _17797_/Q vssd1 vssd1 vccd1 vccd1 _15047_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_115_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16094_ _16096_/A1 _16093_/Y _17725_/C1 vssd1 vssd1 vccd1 vccd1 _18749_/D sky130_fd_sc_hd__a21oi_1
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15045_ _18531_/Q _18530_/Q _17159_/A _15044_/X vssd1 vssd1 vccd1 vccd1 _15045_/X
+ sky130_fd_sc_hd__a211o_1
X_12257_ _16811_/A _12257_/B vssd1 vssd1 vccd1 vccd1 _12257_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ _11201_/X _11207_/X _11622_/C1 vssd1 vssd1 vccd1 vccd1 _11208_/X sky130_fd_sc_hd__a21o_1
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12188_ _17859_/Q _12186_/B _12187_/Y vssd1 vssd1 vccd1 vccd1 _17859_/D sky130_fd_sc_hd__o21a_1
XFILLER_268_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18804_ _19642_/CLK _18804_/D vssd1 vssd1 vccd1 vccd1 _18804_/Q sky130_fd_sc_hd__dfxtp_1
X_11139_ _13487_/S _11139_/B vssd1 vssd1 vccd1 vccd1 _13485_/A sky130_fd_sc_hd__nor2_4
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16996_ _17571_/A _17044_/A2 _16995_/X _17559_/A vssd1 vssd1 vccd1 vccd1 _19334_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_205_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15947_ input8/X input283/X _15947_/S vssd1 vssd1 vccd1 vccd1 _15947_/X sky130_fd_sc_hd__mux2_1
X_18735_ _18738_/CLK _18735_/D vssd1 vssd1 vccd1 vccd1 _18735_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18666_ _18666_/CLK _18666_/D vssd1 vssd1 vccd1 vccd1 _18666_/Q sky130_fd_sc_hd__dfxtp_1
X_15878_ input261/X _15881_/B vssd1 vssd1 vccd1 vccd1 _15878_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_224_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14829_ _12459_/X _14002_/B _14683_/X _18640_/Q vssd1 vssd1 vccd1 vccd1 _14829_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_17617_ _19488_/Q _15093_/B _17556_/A _17205_/B _17556_/X vssd1 vssd1 vccd1 vccd1
+ _17617_/X sky130_fd_sc_hd__a221o_1
X_18597_ _19148_/CLK _18597_/D vssd1 vssd1 vccd1 vccd1 _18597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17548_ _19520_/Q _17547_/B _17546_/X _17547_/Y _17352_/A vssd1 vssd1 vccd1 vccd1
+ _19520_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17479_ _19507_/Q _17547_/B _17477_/X _17478_/Y _17350_/A vssd1 vssd1 vccd1 vccd1
+ _19507_/D sky130_fd_sc_hd__o221a_1
XFILLER_221_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19218_ _19219_/CLK _19218_/D vssd1 vssd1 vccd1 vccd1 _19218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19149_ _19604_/CLK _19149_/D vssd1 vssd1 vccd1 vccd1 _19149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_62_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19594_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_114_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09804_ _19102_/Q _19134_/Q _11609_/S vssd1 vssd1 vccd1 vccd1 _09804_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09735_ _09735_/A _12609_/B vssd1 vssd1 vccd1 vccd1 _09736_/B sky130_fd_sc_hd__or2_4
XFILLER_28_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ _18598_/Q _18169_/Q _09671_/S vssd1 vssd1 vccd1 vccd1 _09666_/X sky130_fd_sc_hd__mux2_1
XFILLER_270_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _18021_/Q _17989_/Q _10721_/S vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10510_ _10506_/X _10507_/X _10668_/S vssd1 vssd1 vccd1 vccd1 _10510_/X sky130_fd_sc_hd__mux2_1
XFILLER_211_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11490_ _18113_/Q _11490_/B vssd1 vssd1 vccd1 vccd1 _11490_/X sky130_fd_sc_hd__or2_2
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10441_ _18465_/Q _18366_/Q _10667_/S vssd1 vssd1 vccd1 vccd1 _10441_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10372_ _10742_/A1 _10359_/X _10360_/X vssd1 vssd1 vccd1 vccd1 _10372_/X sky130_fd_sc_hd__o21a_1
XFILLER_137_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13160_ _18108_/Q _13159_/C _18109_/Q vssd1 vssd1 vccd1 vccd1 _13161_/B sky130_fd_sc_hd__a21oi_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12111_ _17830_/Q _12112_/C _17831_/Q vssd1 vssd1 vccd1 vccd1 _12113_/B sky130_fd_sc_hd__a21oi_1
Xclkbuf_4_10__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_79_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
X_13091_ _12831_/Y _13090_/Y _13314_/S vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__mux2_1
X_12042_ _17896_/Q _12052_/A2 _12041_/X _13100_/A vssd1 vssd1 vccd1 vccd1 _17798_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1702 _09457_/A vssd1 vssd1 vccd1 vccd1 _11480_/C1 sky130_fd_sc_hd__buf_12
Xfanout1713 _08828_/Y vssd1 vssd1 vccd1 vccd1 _16836_/S sky130_fd_sc_hd__buf_8
XFILLER_2_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1724 _16852_/A vssd1 vssd1 vccd1 vccd1 _12488_/A sky130_fd_sc_hd__buf_4
XFILLER_104_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1735 _18339_/Q vssd1 vssd1 vccd1 vccd1 _09651_/S sky130_fd_sc_hd__buf_4
X_16850_ _16967_/S _16850_/B vssd1 vssd1 vccd1 vccd1 _16850_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1746 _18201_/Q vssd1 vssd1 vccd1 vccd1 _08858_/A sky130_fd_sc_hd__buf_4
Xfanout1757 _09553_/A vssd1 vssd1 vccd1 vccd1 _10689_/S sky130_fd_sc_hd__buf_6
X_15801_ _16326_/A _16194_/B vssd1 vssd1 vccd1 vccd1 _15801_/Y sky130_fd_sc_hd__nor2_2
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1768 _10471_/S vssd1 vssd1 vccd1 vccd1 _11327_/S sky130_fd_sc_hd__buf_6
Xfanout770 _17658_/Y vssd1 vssd1 vccd1 vccd1 _17681_/S sky130_fd_sc_hd__buf_6
XFILLER_266_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1779 _12320_/B vssd1 vssd1 vccd1 vccd1 _10589_/S sky130_fd_sc_hd__clkbuf_16
Xfanout781 _16590_/S vssd1 vssd1 vccd1 vccd1 _16585_/S sky130_fd_sc_hd__buf_12
X_16781_ _19281_/Q _16783_/C _16780_/Y vssd1 vssd1 vccd1 vccd1 _19281_/D sky130_fd_sc_hd__a21oi_1
Xfanout792 _16492_/Y vssd1 vssd1 vccd1 vccd1 _16521_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13993_ _14033_/A1 _13217_/X _13992_/X _14029_/C1 vssd1 vssd1 vccd1 vccd1 _17961_/D
+ sky130_fd_sc_hd__o211a_1
X_18520_ _19291_/CLK _18520_/D vssd1 vssd1 vccd1 vccd1 _18520_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15732_ _19452_/Q _15793_/A2 _17208_/A _15731_/Y vssd1 vssd1 vccd1 vccd1 _15732_/Y
+ sky130_fd_sc_hd__o211ai_1
X_12944_ _12942_/X _12943_/X _13130_/A vssd1 vssd1 vccd1 vccd1 _12945_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _19631_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15663_ _18586_/Q _15662_/C _18587_/Q vssd1 vssd1 vccd1 vccd1 _15664_/B sky130_fd_sc_hd__a21oi_1
XFILLER_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _12873_/Y _12874_/X _13089_/A vssd1 vssd1 vccd1 vccd1 _12875_/X sky130_fd_sc_hd__mux2_1
XANTENNA_130 _11814_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _11840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_152 _11872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _18564_/Q _17461_/A2 _17426_/B1 vssd1 vssd1 vccd1 vccd1 _17402_/X sky130_fd_sc_hd__o21a_1
XFILLER_261_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14614_ _16540_/A0 _18421_/Q _14631_/S vssd1 vssd1 vccd1 vccd1 _18421_/D sky130_fd_sc_hd__mux2_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_163 _12461_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ _11826_/A _11826_/B vssd1 vssd1 vccd1 vccd1 _11827_/C sky130_fd_sc_hd__nor2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _19399_/CLK _18382_/D vssd1 vssd1 vccd1 vccd1 _18382_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_174 _13331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15594_ _18583_/Q _15800_/A2 _15586_/X _15593_/X _17376_/A vssd1 vssd1 vccd1 vccd1
+ _18583_/D sky130_fd_sc_hd__o221a_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _13659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_196 _13872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17333_ _19464_/Q _17575_/A _17345_/S vssd1 vssd1 vccd1 vccd1 _17334_/B sky130_fd_sc_hd__mux2_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _18381_/Q _14589_/A2 _14589_/B1 input40/X vssd1 vssd1 vccd1 vccd1 _14546_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _18575_/Q _11759_/A2 _11844_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _11757_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708_ _18648_/Q _18070_/Q _19089_/Q _18993_/Q _11171_/S _11156_/C1 vssd1 vssd1
+ vccd1 vccd1 _10708_/X sky130_fd_sc_hd__mux4_1
X_17264_ _17262_/Y _17263_/X _17261_/A vssd1 vssd1 vccd1 vccd1 _19438_/D sky130_fd_sc_hd__a21oi_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14476_ _18328_/Q _17680_/A0 _14486_/S vssd1 vssd1 vccd1 vccd1 _18328_/D sky130_fd_sc_hd__mux2_1
X_11688_ _18405_/Q _18406_/Q vssd1 vssd1 vccd1 vccd1 _14528_/B sky130_fd_sc_hd__nand2b_4
X_19003_ _19618_/CLK _19003_/D vssd1 vssd1 vccd1 vccd1 _19003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16215_ _17712_/A0 _18831_/Q _16226_/S vssd1 vssd1 vccd1 vccd1 _18831_/D sky130_fd_sc_hd__mux2_1
X_13427_ _13427_/A1 _13425_/X _13952_/B1 vssd1 vssd1 vccd1 vccd1 _13427_/X sky130_fd_sc_hd__a21o_2
X_17195_ _17198_/A _17195_/B vssd1 vssd1 vccd1 vccd1 _19416_/D sky130_fd_sc_hd__nor2_1
X_10639_ _09140_/S _11869_/A _11181_/B1 vssd1 vssd1 vccd1 vccd1 _10639_/X sky130_fd_sc_hd__a21o_1
X_16146_ _18776_/Q _18774_/Q _16145_/X vssd1 vssd1 vccd1 vccd1 _16146_/X sky130_fd_sc_hd__or3b_1
XFILLER_115_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13358_ _13358_/A1 _13357_/X _11446_/B vssd1 vssd1 vccd1 vccd1 _13358_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12309_ _14687_/A _14687_/B _12482_/S vssd1 vssd1 vccd1 vccd1 _14854_/D sky130_fd_sc_hd__and3b_1
XFILLER_170_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16077_ _18741_/Q _16020_/A _16068_/X _16076_/X _14427_/B vssd1 vssd1 vccd1 vccd1
+ _18741_/D sky130_fd_sc_hd__o221a_1
X_13289_ _13289_/A _13289_/B vssd1 vssd1 vccd1 vccd1 _13289_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15028_ _18517_/Q input194/X _15038_/S vssd1 vssd1 vccd1 vccd1 _18517_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput3 coreIndex[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_8
X_16979_ _17217_/B vssd1 vssd1 vccd1 vccd1 _16979_/Y sky130_fd_sc_hd__inv_2
XFILLER_284_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09520_ _10275_/S _09512_/X _09511_/X _08967_/S vssd1 vssd1 vccd1 vccd1 _09520_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18718_ _18772_/CLK _18718_/D vssd1 vssd1 vccd1 vccd1 _18718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_180_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18734_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09451_ _10315_/S _09449_/X _09450_/X _10260_/B1 vssd1 vssd1 vccd1 vccd1 _09451_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_37_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18649_ _19092_/CLK _18649_/D vssd1 vssd1 vccd1 vccd1 _18649_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09382_ _09378_/X _09381_/X _10746_/S vssd1 vssd1 vccd1 vccd1 _09382_/X sky130_fd_sc_hd__mux2_1
XFILLER_212_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput340 _11836_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[15] sky130_fd_sc_hd__buf_4
XFILLER_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput351 _11882_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[25] sky130_fd_sc_hd__buf_4
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput362 _11799_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[6] sky130_fd_sc_hd__buf_4
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput373 _11722_/X vssd1 vssd1 vccd1 vccd1 csb0[1] sky130_fd_sc_hd__buf_4
XFILLER_248_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1009 _16488_/S vssd1 vssd1 vccd1 vccd1 _16490_/S sky130_fd_sc_hd__buf_12
Xoutput384 _11937_/X vssd1 vssd1 vccd1 vccd1 din0[17] sky130_fd_sc_hd__buf_4
Xoutput395 _11947_/X vssd1 vssd1 vccd1 vccd1 din0[27] sky130_fd_sc_hd__buf_4
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ _09716_/X _09717_/X _09718_/S vssd1 vssd1 vccd1 vccd1 _09718_/X sky130_fd_sc_hd__mux2_1
XFILLER_228_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10990_ _18989_/Q _11479_/B vssd1 vssd1 vccd1 vccd1 _10990_/X sky130_fd_sc_hd__or2_1
XFILLER_255_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09649_ input151/X input136/X _09990_/S vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__mux2_8
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12660_ _10159_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _12660_/X sky130_fd_sc_hd__and2b_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11609_/X _11610_/X _11611_/S vssd1 vssd1 vccd1 vccd1 _11611_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12591_ _13462_/A _12585_/X _12590_/Y _13421_/A vssd1 vssd1 vccd1 vccd1 _12591_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_51_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14330_ _18187_/Q _17714_/A0 _14335_/S vssd1 vssd1 vccd1 vccd1 _18187_/D sky130_fd_sc_hd__mux2_1
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11542_ _12638_/A _11669_/B _13697_/A _11540_/X vssd1 vssd1 vccd1 vccd1 _11642_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14261_ _18302_/Q _14261_/A2 _14260_/X _14450_/B vssd1 vssd1 vccd1 vccd1 _18128_/D
+ sky130_fd_sc_hd__o211a_1
X_11473_ _19207_/Q _11482_/A2 _11472_/X _12488_/B vssd1 vssd1 vccd1 vccd1 _11473_/X
+ sky130_fd_sc_hd__a211o_1
X_16000_ _18715_/Q _16002_/A2 _16002_/B1 _18764_/Q _16004_/C1 vssd1 vssd1 vccd1 vccd1
+ _16000_/X sky130_fd_sc_hd__a221o_1
XFILLER_143_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13212_ _19337_/Q _13246_/A2 _13950_/B1 _19465_/Q _13950_/C1 vssd1 vssd1 vccd1 vccd1
+ _13212_/X sky130_fd_sc_hd__a221o_1
X_10424_ _19125_/Q _19157_/Q _10424_/S vssd1 vssd1 vccd1 vccd1 _10424_/X sky130_fd_sc_hd__mux2_1
X_14192_ _18707_/Q _18094_/Q _14200_/S vssd1 vssd1 vccd1 vccd1 _14193_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13143_ _11745_/B _13358_/A1 _13142_/X vssd1 vssd1 vccd1 vccd1 _13143_/Y sky130_fd_sc_hd__o21ai_1
X_10355_ _10200_/S _10353_/X _10354_/X _10356_/C1 vssd1 vssd1 vccd1 vccd1 _10355_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13074_ _17829_/Q _13105_/B _13072_/X _13073_/X _12548_/X vssd1 vssd1 vccd1 vccd1
+ _13074_/X sky130_fd_sc_hd__o221a_2
X_10286_ _11199_/S1 _10280_/X _10283_/X _08904_/A vssd1 vssd1 vccd1 vccd1 _10286_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17951_ _17951_/CLK _17951_/D vssd1 vssd1 vccd1 vccd1 _17951_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1510 _10199_/S vssd1 vssd1 vccd1 vccd1 _10206_/S sky130_fd_sc_hd__buf_6
X_16902_ _16970_/A1 _17934_/Q _16901_/X vssd1 vssd1 vccd1 vccd1 _17587_/A sky130_fd_sc_hd__o21a_4
X_12025_ _17790_/Q _12051_/B vssd1 vssd1 vccd1 vccd1 _12025_/X sky130_fd_sc_hd__or2_1
Xfanout1521 _11503_/S0 vssd1 vssd1 vccd1 vccd1 _10424_/S sky130_fd_sc_hd__buf_6
X_17882_ _19323_/CLK _17882_/D vssd1 vssd1 vccd1 vccd1 _17882_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1532 _10653_/A1 vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__buf_6
XFILLER_250_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1543 _10649_/A1 vssd1 vssd1 vccd1 vccd1 _11606_/S sky130_fd_sc_hd__buf_8
XFILLER_78_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1554 _08899_/Y vssd1 vssd1 vccd1 vccd1 _10280_/S sky130_fd_sc_hd__buf_6
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1565 _08898_/Y vssd1 vssd1 vccd1 vccd1 _11515_/B1 sky130_fd_sc_hd__clkbuf_16
XFILLER_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19621_ _19621_/CLK _19621_/D vssd1 vssd1 vccd1 vccd1 _19621_/Q sky130_fd_sc_hd__dfxtp_1
X_16833_ _16821_/A _17817_/Q _12492_/X vssd1 vssd1 vccd1 vccd1 _17051_/C sky130_fd_sc_hd__a21o_1
XFILLER_65_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1576 fanout1581/X vssd1 vssd1 vccd1 vccd1 _09429_/S sky130_fd_sc_hd__buf_8
XFILLER_254_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1587 _09978_/A1 vssd1 vssd1 vccd1 vccd1 _11199_/S1 sky130_fd_sc_hd__buf_8
Xfanout1598 _08893_/Y vssd1 vssd1 vccd1 vccd1 _08950_/A sky130_fd_sc_hd__buf_6
XFILLER_266_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16764_ _19275_/Q _16767_/C _16764_/B1 vssd1 vssd1 vccd1 vccd1 _16764_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_207_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19552_ _19552_/CLK _19552_/D vssd1 vssd1 vccd1 vccd1 _19552_/Q sky130_fd_sc_hd__dfxtp_1
X_13976_ _14034_/B _13976_/B vssd1 vssd1 vccd1 vccd1 _13976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18503_ _19464_/CLK _18503_/D vssd1 vssd1 vccd1 vccd1 _18503_/Q sky130_fd_sc_hd__dfxtp_1
X_15715_ _15715_/A _15715_/B vssd1 vssd1 vccd1 vccd1 _15715_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12927_ _13028_/C _12927_/B vssd1 vssd1 vccd1 vccd1 _12927_/Y sky130_fd_sc_hd__nor2_1
X_16695_ _19251_/Q _19250_/Q _16695_/C vssd1 vssd1 vccd1 vccd1 _16697_/B sky130_fd_sc_hd__and3_1
X_19483_ _19483_/CLK _19483_/D vssd1 vssd1 vccd1 vccd1 _19483_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18434_ _19596_/CLK _18434_/D vssd1 vssd1 vccd1 vccd1 _18434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15646_ _18586_/Q _15662_/C vssd1 vssd1 vccd1 vccd1 _15646_/Y sky130_fd_sc_hd__xnor2_1
X_12858_ _19298_/Q _12583_/Y _12584_/Y input3/X _12857_/X vssd1 vssd1 vccd1 vccd1
+ _12858_/X sky130_fd_sc_hd__a221o_4
XFILLER_179_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ _19641_/CLK _18365_/D vssd1 vssd1 vccd1 vccd1 _18365_/Q sky130_fd_sc_hd__dfxtp_1
X_11809_ _11820_/A _11808_/X _11807_/Y vssd1 vssd1 vccd1 vccd1 _11810_/C sky130_fd_sc_hd__a21oi_4
X_15577_ _15787_/A _15639_/A vssd1 vssd1 vccd1 vccd1 _15577_/X sky130_fd_sc_hd__and2_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12868_/B _12789_/B vssd1 vssd1 vccd1 vccd1 _12790_/A sky130_fd_sc_hd__nor2_1
XFILLER_221_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17316_ _17316_/A _17316_/B vssd1 vssd1 vccd1 vccd1 _17337_/S sky130_fd_sc_hd__nor2_8
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14528_ _14528_/A _14528_/B vssd1 vssd1 vccd1 vccd1 _14528_/X sky130_fd_sc_hd__or2_1
X_18296_ _19453_/CLK _18296_/D vssd1 vssd1 vccd1 vccd1 _18296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17247_ _19433_/Q _17310_/B vssd1 vssd1 vccd1 vccd1 _17247_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14459_ _18311_/Q _17663_/A0 _14483_/S vssd1 vssd1 vccd1 vccd1 _18311_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17178_ _17208_/A _17178_/B vssd1 vssd1 vccd1 vccd1 _17488_/A sky130_fd_sc_hd__nand2_1
XFILLER_183_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16129_ _18767_/Q _16139_/B vssd1 vssd1 vccd1 vccd1 _16129_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08951_ _11198_/S _14350_/A vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__xnor2_1
XFILLER_170_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08882_ _10027_/A _08882_/B vssd1 vssd1 vccd1 vccd1 _08882_/Y sky130_fd_sc_hd__nand2_2
XFILLER_96_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09503_ _19624_/Q _18913_/Q _09952_/S vssd1 vssd1 vccd1 vccd1 _09503_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09434_ _17927_/Q _08947_/X _09433_/X vssd1 vssd1 vccd1 vccd1 _09434_/X sky130_fd_sc_hd__a21o_2
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ _09643_/A _11804_/A vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__and2_2
XFILLER_200_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09296_ _09292_/X _09295_/X _10746_/S vssd1 vssd1 vccd1 vccd1 _09296_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_30 _17205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 _11812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_52 _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_63 _13917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_74 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_85 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_96 _13515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ _18266_/Q _18841_/Q _10141_/S vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10071_ _09736_/B _10070_/A _10070_/B _09734_/Y vssd1 vssd1 vccd1 vccd1 _11739_/B
+ sky130_fd_sc_hd__a31o_4
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13830_ _13928_/A1 _13819_/X _13821_/Y _13829_/Y vssd1 vssd1 vccd1 vccd1 _14028_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_275_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ _13761_/A _13761_/B vssd1 vssd1 vccd1 vccd1 _13761_/X sky130_fd_sc_hd__or2_1
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10973_ _10971_/X _10972_/X _11361_/S vssd1 vssd1 vccd1 vccd1 _10973_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15500_ _18579_/Q _15447_/B _15492_/X _15499_/X _17350_/A vssd1 vssd1 vccd1 vccd1
+ _18579_/D sky130_fd_sc_hd__o221a_1
XFILLER_188_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12712_ _12609_/B _12653_/B _12712_/S vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _17679_/A0 _19087_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _19087_/D sky130_fd_sc_hd__mux2_1
X_13692_ _13929_/A1 _13691_/X _13679_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_243_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15431_ _15432_/A _15432_/B vssd1 vssd1 vccd1 vccd1 _15431_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12643_ _13665_/A _12643_/B vssd1 vssd1 vccd1 vccd1 _12643_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18150_ _19635_/CLK _18150_/D vssd1 vssd1 vccd1 vccd1 _18150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15362_ _15289_/A _15289_/B _15262_/A _15262_/B vssd1 vssd1 vccd1 vccd1 _15362_/X
+ sky130_fd_sc_hd__a211o_1
X_12574_ _12582_/A _12576_/B vssd1 vssd1 vccd1 vccd1 _12918_/S sky130_fd_sc_hd__nor2_4
XFILLER_30_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17101_ _19384_/Q _17107_/B vssd1 vssd1 vccd1 vccd1 _17101_/X sky130_fd_sc_hd__or2_1
XFILLER_196_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14313_ _18170_/Q _17697_/A0 _14335_/S vssd1 vssd1 vccd1 vccd1 _18170_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18081_ _18746_/CLK _18081_/D vssd1 vssd1 vccd1 vccd1 _18081_/Q sky130_fd_sc_hd__dfxtp_1
X_11525_ _09145_/A _10080_/B _13267_/A vssd1 vssd1 vccd1 vccd1 _11681_/B sky130_fd_sc_hd__o21ba_4
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15293_ _15365_/B _15293_/B vssd1 vssd1 vccd1 vccd1 _15293_/X sky130_fd_sc_hd__xor2_1
XFILLER_157_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17032_ _17193_/B _17032_/A2 _17031_/X _17366_/A vssd1 vssd1 vccd1 vccd1 _19352_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14244_ _18120_/Q _14244_/B vssd1 vssd1 vccd1 vccd1 _14244_/X sky130_fd_sc_hd__or2_1
X_11456_ _10403_/S _11455_/X _11454_/X _09135_/S vssd1 vssd1 vccd1 vccd1 _11456_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ _11458_/A1 _19157_/Q _11379_/S _19125_/Q vssd1 vssd1 vccd1 vccd1 _10407_/X
+ sky130_fd_sc_hd__o22a_1
X_14175_ _16968_/A _14175_/B vssd1 vssd1 vccd1 vccd1 _18085_/D sky130_fd_sc_hd__and2_1
XFILLER_139_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11387_ _11464_/C1 _11386_/X _11385_/X _11478_/S vssd1 vssd1 vccd1 vccd1 _11387_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13126_ _13126_/A _13126_/B vssd1 vssd1 vccd1 vccd1 _13127_/B sky130_fd_sc_hd__nand2_1
X_10338_ _10338_/A1 _10337_/X _11459_/B1 vssd1 vssd1 vccd1 vccd1 _10338_/X sky130_fd_sc_hd__o21a_1
XFILLER_152_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18983_ _19079_/CLK _18983_/D vssd1 vssd1 vccd1 vccd1 _18983_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19327_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _18749_/CLK _17934_/D vssd1 vssd1 vccd1 vccd1 _17934_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _15330_/A _13056_/X _13237_/B1 vssd1 vssd1 vccd1 vccd1 _13057_/Y sky130_fd_sc_hd__o21ai_1
X_10269_ _10180_/A _10247_/X _10255_/Y _10261_/Y _10268_/Y vssd1 vssd1 vccd1 vccd1
+ _10269_/X sky130_fd_sc_hd__a32o_2
XFILLER_79_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1340 _09096_/Y vssd1 vssd1 vccd1 vccd1 _10004_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ _17775_/Q _17709_/A0 _12022_/S vssd1 vssd1 vccd1 vccd1 _17775_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1351 _09919_/C1 vssd1 vssd1 vccd1 vccd1 _10338_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_239_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17865_ _17865_/CLK _17865_/D vssd1 vssd1 vccd1 vccd1 _17865_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1362 _09093_/Y vssd1 vssd1 vccd1 vccd1 _11167_/B sky130_fd_sc_hd__buf_8
XFILLER_94_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1373 _10467_/S vssd1 vssd1 vccd1 vccd1 _10613_/S sky130_fd_sc_hd__buf_6
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1384 fanout1386/X vssd1 vssd1 vccd1 vccd1 _11226_/S sky130_fd_sc_hd__buf_6
X_19604_ _19604_/CLK _19604_/D vssd1 vssd1 vccd1 vccd1 _19604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16816_ _16964_/A _16816_/B _16816_/C vssd1 vssd1 vccd1 vccd1 _19294_/D sky130_fd_sc_hd__and3_1
Xfanout1395 fanout1407/X vssd1 vssd1 vccd1 vccd1 _10320_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17796_ _19650_/CLK _17796_/D vssd1 vssd1 vccd1 vccd1 _17796_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19535_ _19552_/CLK _19535_/D vssd1 vssd1 vccd1 vccd1 _19535_/Q sky130_fd_sc_hd__dfxtp_1
X_16747_ _16752_/A _16747_/B _16751_/C vssd1 vssd1 vccd1 vccd1 _19268_/D sky130_fd_sc_hd__nor3_1
X_13959_ _12656_/A _13908_/B _12660_/X _12656_/B vssd1 vssd1 vccd1 vccd1 _13959_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_235_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16678_ _16776_/A _16688_/C vssd1 vssd1 vccd1 vccd1 _16678_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19466_ _19466_/CLK _19466_/D vssd1 vssd1 vccd1 vccd1 _19466_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_222_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18417_ _19564_/CLK _18417_/D vssd1 vssd1 vccd1 vccd1 _18417_/Q sky130_fd_sc_hd__dfxtp_1
X_15629_ _19479_/Q _19413_/Q vssd1 vssd1 vccd1 vccd1 _15630_/B sky130_fd_sc_hd__or2_1
X_19397_ _19466_/CLK _19397_/D vssd1 vssd1 vccd1 vccd1 _19397_/Q sky130_fd_sc_hd__dfxtp_2
X_09150_ _09908_/A1 _09236_/A _09149_/X _09908_/B1 _18391_/Q vssd1 vssd1 vccd1 vccd1
+ _09150_/X sky130_fd_sc_hd__o32a_1
XFILLER_194_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18348_ _19213_/CLK _18348_/D vssd1 vssd1 vccd1 vccd1 _18348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18279_ _18279_/CLK _18279_/D vssd1 vssd1 vccd1 vccd1 _18279_/Q sky130_fd_sc_hd__dfxtp_1
X_09081_ _12445_/A _13294_/A vssd1 vssd1 vccd1 vccd1 _09697_/B sky130_fd_sc_hd__nand2_4
XFILLER_175_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput50 dout0[16] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_2
XFILLER_238_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput61 dout0[26] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
Xinput72 dout0[36] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput83 dout0[46] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_2
Xinput94 dout0[56] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09983_ _09984_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _14141_/A sky130_fd_sc_hd__xnor2_4
XFILLER_254_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08934_ _17819_/Q _17818_/Q _17817_/Q _17816_/Q vssd1 vssd1 vccd1 vccd1 _08935_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_258_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08865_ _18080_/Q _17887_/Q vssd1 vssd1 vccd1 vccd1 _08865_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_111_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09417_ _10300_/S _09414_/X _09416_/X vssd1 vssd1 vccd1 vccd1 _09417_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_241_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09348_ _10262_/A1 _19626_/Q _18915_/Q _10099_/S vssd1 vssd1 vccd1 vccd1 _09348_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _17917_/Q _09643_/A vssd1 vssd1 vccd1 vccd1 _09279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11310_ _11311_/C1 _11309_/X _11308_/X _10930_/S vssd1 vssd1 vccd1 vccd1 _11310_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_154_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12290_ _12486_/B _12457_/B vssd1 vssd1 vccd1 vccd1 _12292_/C sky130_fd_sc_hd__or2_2
XFILLER_154_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11241_ _19050_/Q _19018_/Q _11247_/S vssd1 vssd1 vccd1 vccd1 _11241_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11172_ _11172_/A1 _18149_/Q _18795_/Q _11171_/S vssd1 vssd1 vccd1 vccd1 _11172_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ _18337_/Q _17788_/Q _10206_/S vssd1 vssd1 vccd1 vccd1 _10123_/X sky130_fd_sc_hd__mux2_1
X_15980_ _18705_/Q _15953_/B _16004_/B1 _18754_/Q _16004_/C1 vssd1 vssd1 vccd1 vccd1
+ _15980_/X sky130_fd_sc_hd__a221o_1
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10054_ _19067_/Q _18971_/Q _10054_/S vssd1 vssd1 vccd1 vccd1 _10054_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14931_ _17814_/Q _15002_/B vssd1 vssd1 vccd1 vccd1 _14931_/X sky130_fd_sc_hd__or2_1
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17650_ _17683_/A0 _19578_/Q _17657_/S vssd1 vssd1 vccd1 vccd1 _19578_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14862_ _15003_/A1 _13505_/Y _15003_/B1 _18643_/Q _15003_/C1 vssd1 vssd1 vccd1 vccd1
+ _14862_/X sky130_fd_sc_hd__a221o_1
XFILLER_275_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _17668_/A0 _19204_/Q _16622_/S vssd1 vssd1 vccd1 vccd1 _19204_/D sky130_fd_sc_hd__mux2_1
X_13813_ _13861_/A _14152_/A _13892_/B1 vssd1 vssd1 vccd1 vccd1 _13813_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17581_ _17581_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17581_/X sky130_fd_sc_hd__or2_1
XFILLER_251_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14793_ _14865_/A1 _14792_/X _14865_/B1 vssd1 vssd1 vccd1 vccd1 _14793_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19320_ _19320_/CLK _19320_/D vssd1 vssd1 vccd1 vccd1 _19320_/Q sky130_fd_sc_hd__dfxtp_1
X_16532_ _16532_/A0 _19137_/Q _16548_/S vssd1 vssd1 vccd1 vccd1 _19137_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13744_ _17848_/Q _13744_/A2 _13744_/B1 _17880_/Q vssd1 vssd1 vccd1 vccd1 _13744_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10956_ _11355_/A1 _10955_/X _11608_/C1 vssd1 vssd1 vccd1 vccd1 _10956_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19251_ _19261_/CLK _19251_/D vssd1 vssd1 vccd1 vccd1 _19251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16463_ _16529_/A0 _19070_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _19070_/D sky130_fd_sc_hd__mux2_1
X_13675_ _13739_/A _13675_/B vssd1 vssd1 vccd1 vccd1 _13675_/Y sky130_fd_sc_hd__nand2_2
XFILLER_232_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10887_ _10887_/A _10887_/B vssd1 vssd1 vccd1 vccd1 _10887_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18202_ _19231_/CLK _18202_/D vssd1 vssd1 vccd1 vccd1 _18202_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15414_ _15465_/C _15414_/B vssd1 vssd1 vccd1 vccd1 _15416_/B sky130_fd_sc_hd__nor2_1
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19182_ _19637_/CLK _19182_/D vssd1 vssd1 vccd1 vccd1 _19182_/Q sky130_fd_sc_hd__dfxtp_1
X_12626_ _12626_/A _12626_/B _13351_/A _13311_/A vssd1 vssd1 vccd1 vccd1 _12626_/X
+ sky130_fd_sc_hd__or4_1
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16394_ _17692_/A0 _19003_/Q _16425_/S vssd1 vssd1 vccd1 vccd1 _19003_/D sky130_fd_sc_hd__mux2_1
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18133_ _19099_/CLK _18133_/D vssd1 vssd1 vccd1 vccd1 _18133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15345_ _19467_/Q _19401_/Q vssd1 vssd1 vccd1 vccd1 _15347_/A sky130_fd_sc_hd__xnor2_1
XFILLER_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _12768_/B _12561_/B vssd1 vssd1 vccd1 vccd1 _12557_/X sky130_fd_sc_hd__or2_1
X_11508_ _11428_/A _11507_/X _11508_/B1 vssd1 vssd1 vccd1 vccd1 _11509_/B sky130_fd_sc_hd__a21o_1
XFILLER_144_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18064_ _19197_/CLK _18064_/D vssd1 vssd1 vccd1 vccd1 _18064_/Q sky130_fd_sc_hd__dfxtp_1
X_15276_ _19464_/Q _19398_/Q vssd1 vssd1 vccd1 vccd1 _15277_/B sky130_fd_sc_hd__nand2_2
X_12488_ _12488_/A _12488_/B vssd1 vssd1 vccd1 vccd1 _12488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17015_ _19344_/Q _17045_/B vssd1 vssd1 vccd1 vccd1 _17015_/X sky130_fd_sc_hd__or2_1
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14227_ _18285_/Q _14267_/A2 _14226_/X _14452_/B vssd1 vssd1 vccd1 vccd1 _18111_/D
+ sky130_fd_sc_hd__o211a_1
X_11439_ _11053_/A _11418_/Y _11424_/Y _11431_/Y _11438_/X vssd1 vssd1 vccd1 vccd1
+ _11439_/X sky130_fd_sc_hd__o32a_4
XFILLER_208_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14158_ _14158_/A _14158_/B _14158_/C vssd1 vssd1 vccd1 vccd1 _15328_/C sky130_fd_sc_hd__or3_4
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13109_ _19399_/Q _12570_/A _13244_/B1 vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__a21o_1
X_14089_ _17672_/A0 _18029_/Q _14104_/S vssd1 vssd1 vccd1 vccd1 _18029_/D sky130_fd_sc_hd__mux2_1
X_18966_ _19596_/CLK _18966_/D vssd1 vssd1 vccd1 vccd1 _18966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17917_ _18881_/CLK _17917_/D vssd1 vssd1 vccd1 vccd1 _17917_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18897_ _19601_/CLK _18897_/D vssd1 vssd1 vccd1 vccd1 _18897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1170 _15851_/Y vssd1 vssd1 vccd1 vccd1 _15948_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_239_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1181 _15304_/A1 vssd1 vssd1 vccd1 vccd1 _15259_/B sky130_fd_sc_hd__clkbuf_8
Xfanout1192 _16002_/B1 vssd1 vssd1 vccd1 vccd1 _16004_/B1 sky130_fd_sc_hd__buf_4
X_17848_ _19324_/CLK _17848_/D vssd1 vssd1 vccd1 vccd1 _17848_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17975_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17779_ _19575_/CLK _17779_/D vssd1 vssd1 vccd1 vccd1 _17779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19518_ _19519_/CLK _19518_/D vssd1 vssd1 vccd1 vccd1 _19518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19586_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_241_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19449_ _19484_/CLK _19449_/D vssd1 vssd1 vccd1 vccd1 _19449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09202_ _10297_/A1 _09199_/X _09200_/X vssd1 vssd1 vccd1 vccd1 _09203_/B sky130_fd_sc_hd__o21ai_1
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09133_ _09130_/X _09132_/X _09135_/S vssd1 vssd1 vccd1 vccd1 _09133_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09064_ _12756_/A _12264_/A vssd1 vssd1 vccd1 vccd1 _12665_/B sky130_fd_sc_hd__or2_2
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09966_ _18533_/Q _18408_/Q _09966_/S vssd1 vssd1 vccd1 vccd1 _09966_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08917_ _08816_/A _17801_/Q vssd1 vssd1 vccd1 vccd1 _14488_/B sky130_fd_sc_hd__nand2b_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _09898_/A _12602_/B vssd1 vssd1 vccd1 vccd1 _09897_/Y sky130_fd_sc_hd__nor2_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _08896_/A vssd1 vssd1 vccd1 vccd1 _08848_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_217_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_504 _10027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_515 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_526 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_537 input231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810_ _18257_/Q _18832_/Q _11598_/S vssd1 vssd1 vccd1 vccd1 _10810_/X sky130_fd_sc_hd__mux2_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_548 _12320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11790_ _15081_/A _11790_/B _11790_/C _11790_/D vssd1 vssd1 vccd1 vccd1 wire989/A
+ sky130_fd_sc_hd__nor4_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10741_ _10373_/S _10736_/X _10740_/X _08895_/A vssd1 vssd1 vccd1 vccd1 _10741_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13460_ _12454_/X _14006_/B _13446_/Y vssd1 vssd1 vccd1 vccd1 _13462_/B sky130_fd_sc_hd__o21ai_1
XFILLER_230_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10672_ _11279_/B1 _10655_/X _10670_/X _10671_/Y vssd1 vssd1 vccd1 vccd1 _10672_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_201_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12411_ _12429_/A1 _09232_/A _09320_/X _12417_/B1 _18397_/Q vssd1 vssd1 vccd1 vccd1
+ _12412_/B sky130_fd_sc_hd__o32ai_4
X_13391_ _13136_/S _12828_/X _13197_/B1 vssd1 vssd1 vccd1 vccd1 _13391_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_166_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15130_ _15130_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15130_/X sky130_fd_sc_hd__and2_1
XFILLER_127_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12342_ _18374_/Q _12432_/B1 _09907_/Y _08858_/A vssd1 vssd1 vccd1 vccd1 _12343_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15061_ _18545_/Q _17672_/A0 _15078_/S vssd1 vssd1 vccd1 vccd1 _18545_/D sky130_fd_sc_hd__mux2_1
XFILLER_182_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12273_ _18775_/Q _18774_/Q _18776_/Q vssd1 vssd1 vccd1 vccd1 _15835_/C sky130_fd_sc_hd__or3b_4
XFILLER_175_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14012_ _14020_/B _14012_/B vssd1 vssd1 vccd1 vccd1 _14012_/Y sky130_fd_sc_hd__nand2_1
X_11224_ _18986_/Q _11224_/B vssd1 vssd1 vccd1 vccd1 _11224_/X sky130_fd_sc_hd__or2_1
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18820_ _19206_/CLK _18820_/D vssd1 vssd1 vccd1 vccd1 _18820_/Q sky130_fd_sc_hd__dfxtp_1
X_11155_ _11156_/C1 _11154_/X _11153_/X _11161_/S vssd1 vssd1 vccd1 vccd1 _11155_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10106_ _18562_/Q _18437_/Q _18046_/Q _18014_/Q _10090_/S _11001_/C1 vssd1 vssd1
+ vccd1 vccd1 _10106_/X sky130_fd_sc_hd__mux4_1
X_18751_ _18776_/CLK _18751_/D vssd1 vssd1 vccd1 vccd1 _18751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15963_ _18697_/Q _15977_/A2 _15962_/X _16892_/A vssd1 vssd1 vccd1 vccd1 _18697_/D
+ sky130_fd_sc_hd__o211a_1
X_11086_ _11251_/S _19180_/Q _11094_/S vssd1 vssd1 vccd1 vccd1 _11086_/X sky130_fd_sc_hd__and3_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput240 localMemory_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input240/X sky130_fd_sc_hd__buf_8
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput251 localMemory_wb_stb_i vssd1 vssd1 vccd1 vccd1 _15013_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17702_ _17702_/A0 _19628_/Q _17722_/S vssd1 vssd1 vccd1 vccd1 _19628_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput262 manufacturerID[8] vssd1 vssd1 vccd1 vccd1 _15881_/A sky130_fd_sc_hd__buf_4
XFILLER_209_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14914_ _18123_/Q _14801_/B _14852_/X _14913_/X vssd1 vssd1 vccd1 vccd1 _14914_/X
+ sky130_fd_sc_hd__o211a_1
X_10037_ _10033_/X _10036_/X _10589_/S vssd1 vssd1 vccd1 vccd1 _10037_/X sky130_fd_sc_hd__mux2_1
Xinput273 partID[3] vssd1 vssd1 vccd1 vccd1 _15899_/A sky130_fd_sc_hd__clkbuf_2
X_18682_ _18683_/CLK _18682_/D vssd1 vssd1 vccd1 vccd1 _18682_/Q sky130_fd_sc_hd__dfxtp_1
X_15894_ _18673_/Q _15906_/A2 _15903_/B1 _15893_/X vssd1 vssd1 vccd1 vccd1 _15894_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput284 wb_rst_i vssd1 vssd1 vccd1 vccd1 input284/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _17666_/A0 _19561_/Q _17654_/S vssd1 vssd1 vccd1 vccd1 _19561_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14845_ _14845_/A vssd1 vssd1 vccd1 vccd1 _14845_/Y sky130_fd_sc_hd__clkinv_4
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17564_ _19524_/Q _17561_/B _17588_/B1 _17563_/X vssd1 vssd1 vccd1 vccd1 _19524_/D
+ sky130_fd_sc_hd__o211a_1
X_14776_ _14696_/A _18270_/Q _14775_/Y _14846_/B1 vssd1 vssd1 vccd1 vccd1 _14776_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_223_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11988_ _14074_/C _14272_/B vssd1 vssd1 vccd1 vccd1 _14351_/A sky130_fd_sc_hd__or2_4
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19303_ _19326_/CLK _19303_/D vssd1 vssd1 vccd1 vccd1 _19303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13727_ _13727_/A _13727_/B vssd1 vssd1 vccd1 vccd1 _14148_/B sky130_fd_sc_hd__xnor2_2
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16515_ _16548_/A0 _19121_/Q _16515_/S vssd1 vssd1 vccd1 vccd1 _19121_/D sky130_fd_sc_hd__mux2_1
XFILLER_205_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10939_ _10930_/S _10938_/X _11328_/S vssd1 vssd1 vccd1 vccd1 _10939_/X sky130_fd_sc_hd__a21o_1
XFILLER_260_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17495_ _13622_/B _17520_/A2 _17543_/B1 _17811_/Q _17550_/A vssd1 vssd1 vccd1 vccd1
+ _17495_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19234_ _19268_/CLK _19234_/D vssd1 vssd1 vccd1 vccd1 _19234_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_220_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13658_ _19318_/Q _13174_/A _13722_/B1 _13651_/X _13657_/X vssd1 vssd1 vccd1 vccd1
+ _13658_/Y sky130_fd_sc_hd__a2111oi_2
X_16446_ _19054_/Q _16611_/A0 _16453_/S vssd1 vssd1 vccd1 vccd1 _19054_/D sky130_fd_sc_hd__mux2_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _12609_/A _12609_/B vssd1 vssd1 vccd1 vccd1 _12610_/B sky130_fd_sc_hd__nand2_1
X_16377_ _16543_/A0 _18988_/Q _16391_/S vssd1 vssd1 vccd1 vccd1 _18988_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19165_ _19197_/CLK _19165_/D vssd1 vssd1 vccd1 vccd1 _19165_/Q sky130_fd_sc_hd__dfxtp_1
X_13589_ _19444_/Q _13949_/A2 _13587_/X _13588_/X _13949_/C1 vssd1 vssd1 vccd1 vccd1
+ _13589_/X sky130_fd_sc_hd__o221a_1
XFILLER_191_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18116_ _19450_/CLK _18116_/D vssd1 vssd1 vccd1 vccd1 _18116_/Q sky130_fd_sc_hd__dfxtp_4
X_15328_ _17895_/Q _15328_/B _15328_/C vssd1 vssd1 vccd1 vccd1 _15328_/X sky130_fd_sc_hd__and3_1
XFILLER_118_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19096_ _19615_/CLK _19096_/D vssd1 vssd1 vccd1 vccd1 _19096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_134_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19458_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18047_ _19134_/CLK _18047_/D vssd1 vssd1 vccd1 vccd1 _18047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15259_ _15259_/A _15259_/B vssd1 vssd1 vccd1 vccd1 _15259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09820_ _11217_/A _09027_/A _09150_/X _10085_/A vssd1 vssd1 vccd1 vccd1 _09821_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_87_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09751_ _19038_/Q _09770_/S vssd1 vssd1 vccd1 vccd1 _09751_/X sky130_fd_sc_hd__or2_1
X_18949_ _19564_/CLK _18949_/D vssd1 vssd1 vccd1 vccd1 _18949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09682_ _09680_/X _09681_/X _10264_/S vssd1 vssd1 vccd1 vccd1 _09683_/B sky130_fd_sc_hd__mux2_1
XFILLER_239_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09116_ _12408_/A _09114_/X _09115_/X _09264_/S _09112_/X vssd1 vssd1 vccd1 vccd1
+ _09116_/X sky130_fd_sc_hd__o311a_1
XFILLER_136_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09047_ _18384_/Q _11692_/A1 _09331_/A _09046_/Y vssd1 vssd1 vccd1 vccd1 _09047_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1906 input284/X vssd1 vssd1 vccd1 vccd1 _14487_/A sky130_fd_sc_hd__buf_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout930 _15083_/Y vssd1 vssd1 vccd1 vccd1 _17475_/B1 sky130_fd_sc_hd__buf_2
Xfanout941 _14672_/X vssd1 vssd1 vccd1 vccd1 _14973_/C1 sky130_fd_sc_hd__clkbuf_4
X_09949_ _19036_/Q _19004_/Q _09973_/S vssd1 vssd1 vccd1 vccd1 _09949_/X sky130_fd_sc_hd__mux2_1
Xfanout952 _14632_/Y vssd1 vssd1 vccd1 vccd1 _14648_/S sky130_fd_sc_hd__clkbuf_16
Xfanout963 _14137_/S vssd1 vssd1 vccd1 vccd1 _14139_/S sky130_fd_sc_hd__clkbuf_16
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout974 _13527_/B1 vssd1 vssd1 vccd1 vccd1 _13747_/B2 sky130_fd_sc_hd__buf_6
XFILLER_219_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout985 _12450_/Y vssd1 vssd1 vccd1 vccd1 _13808_/C1 sky130_fd_sc_hd__buf_6
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout996 _16617_/A0 vssd1 vssd1 vccd1 vccd1 _17717_/A0 sky130_fd_sc_hd__clkbuf_4
X_12960_ _09780_/X _13292_/A2 _12959_/X _13256_/B1 _17923_/Q vssd1 vssd1 vccd1 vccd1
+ _12961_/B sky130_fd_sc_hd__a32o_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _18565_/Q _11663_/A _11706_/B _12956_/A vssd1 vssd1 vccd1 vccd1 _11911_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_273_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12739_/S _12889_/X _12890_/X vssd1 vssd1 vccd1 vccd1 _12891_/X sky130_fd_sc_hd__a21o_1
XFILLER_46_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 _18101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _16490_/A0 _18437_/Q _14630_/S vssd1 vssd1 vccd1 vccd1 _18437_/D sky130_fd_sc_hd__mux2_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 _18115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11842_ _11859_/B _11786_/Y _11808_/X _14141_/B vssd1 vssd1 vccd1 vccd1 _11842_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 _18107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_334 _16291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_345 _09137_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_356 _12461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 _12053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _18389_/Q _14591_/A2 _14591_/B1 input17/X vssd1 vssd1 vccd1 vccd1 _14562_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_378 _14899_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11865_/A _12265_/B _11816_/A vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__a21oi_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_389 _17591_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _17698_/A0 _18913_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _18913_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13512_ _13904_/A _13512_/B vssd1 vssd1 vccd1 vccd1 _13512_/X sky130_fd_sc_hd__or2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17280_ _19444_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17280_/Y sky130_fd_sc_hd__nand2_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _19121_/Q _19153_/Q _10726_/S vssd1 vssd1 vccd1 vccd1 _10724_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _17661_/A0 _18342_/Q _14521_/S vssd1 vssd1 vccd1 vccd1 _18342_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ _17662_/A0 _18846_/Q _16245_/S vssd1 vssd1 vccd1 vccd1 _18846_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13443_ _13937_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _13443_/X sky130_fd_sc_hd__or2_1
XFILLER_186_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10655_ _11131_/A _10649_/X _10652_/X _10654_/X vssd1 vssd1 vccd1 vccd1 _10655_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16162_ _16592_/A0 _18779_/Q _16165_/S vssd1 vssd1 vccd1 vccd1 _18779_/D sky130_fd_sc_hd__mux2_1
XFILLER_103_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13374_ _19438_/Q _12582_/X _13373_/X vssd1 vssd1 vccd1 vccd1 _13374_/X sky130_fd_sc_hd__o21a_2
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10586_ _18867_/Q _18899_/Q _10656_/S vssd1 vssd1 vccd1 vccd1 _10586_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15113_ _15330_/A _15124_/C vssd1 vssd1 vccd1 vccd1 _15113_/Y sky130_fd_sc_hd__nand2_4
X_12325_ _08943_/Y _12324_/Y _08940_/X vssd1 vssd1 vccd1 vccd1 _12325_/X sky130_fd_sc_hd__a21o_1
XFILLER_86_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16093_ _18749_/Q _16093_/B vssd1 vssd1 vccd1 vccd1 _16093_/Y sky130_fd_sc_hd__nand2_1
XFILLER_182_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15044_ input252/X _15014_/C _15014_/B vssd1 vssd1 vccd1 vccd1 _15044_/X sky130_fd_sc_hd__o21ba_1
X_12256_ _17885_/Q _12256_/B vssd1 vssd1 vccd1 vccd1 _12257_/B sky130_fd_sc_hd__and2_1
XFILLER_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_11207_ _10719_/S _11202_/X _11206_/X vssd1 vssd1 vccd1 vccd1 _11207_/X sky130_fd_sc_hd__a21o_1
XFILLER_122_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12187_ _12187_/A _12192_/C vssd1 vssd1 vccd1 vccd1 _12187_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18803_ _19642_/CLK _18803_/D vssd1 vssd1 vccd1 vccd1 _18803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11138_ _11138_/A _11138_/B vssd1 vssd1 vccd1 vccd1 _11139_/B sky130_fd_sc_hd__nor2_2
XFILLER_268_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16995_ _19334_/Q _17043_/B vssd1 vssd1 vccd1 vccd1 _16995_/X sky130_fd_sc_hd__or2_1
XFILLER_95_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18734_ _18734_/CLK _18734_/D vssd1 vssd1 vccd1 vccd1 _18734_/Q sky130_fd_sc_hd__dfxtp_4
X_15946_ _18691_/Q _15946_/A2 _15945_/X _15946_/C1 vssd1 vssd1 vccd1 vccd1 _18691_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ _19084_/Q _11070_/S _11068_/X _11559_/S1 vssd1 vssd1 vccd1 vccd1 _11069_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18665_ _18666_/CLK _18665_/D vssd1 vssd1 vccd1 vccd1 _18665_/Q sky130_fd_sc_hd__dfxtp_1
X_15877_ _18668_/Q _15949_/A2 _15875_/X _15876_/X _15904_/C1 vssd1 vssd1 vccd1 vccd1
+ _18668_/D sky130_fd_sc_hd__o221a_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17616_ _19549_/Q _17624_/A2 _17615_/X _17592_/B vssd1 vssd1 vccd1 vccd1 _19549_/D
+ sky130_fd_sc_hd__o211a_1
X_14828_ _18484_/Q _15001_/A2 _14827_/Y _12249_/A vssd1 vssd1 vccd1 vccd1 _18484_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18596_ _19588_/CLK _18596_/D vssd1 vssd1 vccd1 vccd1 _18596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17547_ _17547_/A _17547_/B vssd1 vssd1 vccd1 vccd1 _17547_/Y sky130_fd_sc_hd__nand2_1
X_14759_ _17797_/Q _14911_/B vssd1 vssd1 vccd1 vccd1 _14759_/X sky130_fd_sc_hd__or2_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17478_ _17478_/A _17547_/B vssd1 vssd1 vccd1 vccd1 _17478_/Y sky130_fd_sc_hd__nand2_1
X_19217_ _19623_/CLK _19217_/D vssd1 vssd1 vccd1 vccd1 _19217_/Q sky130_fd_sc_hd__dfxtp_1
X_16429_ _19037_/Q _09825_/X _16454_/S vssd1 vssd1 vccd1 vccd1 _19037_/D sky130_fd_sc_hd__mux2_1
X_19148_ _19148_/CLK _19148_/D vssd1 vssd1 vccd1 vccd1 _19148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19079_ _19079_/CLK _19079_/D vssd1 vssd1 vccd1 vccd1 _19079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09803_ _18051_/Q _10816_/A2 _09802_/X _11282_/A vssd1 vssd1 vccd1 vccd1 _09803_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09734_ _12999_/S vssd1 vssd1 vccd1 vccd1 _09734_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_31_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19147_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09665_ _11481_/A _09663_/X _09664_/X vssd1 vssd1 vccd1 vccd1 _09665_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_27_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09596_ _10366_/A1 _19559_/Q _10717_/S _19591_/Q _10371_/S vssd1 vssd1 vccd1 vccd1
+ _09596_/X sky130_fd_sc_hd__o221a_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _10436_/X _10439_/X _11601_/A vssd1 vssd1 vccd1 vccd1 _10440_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _10369_/X _10370_/X _10371_/S vssd1 vssd1 vccd1 vccd1 _10371_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12110_ _17830_/Q _12112_/C _12109_/Y vssd1 vssd1 vccd1 vccd1 _17830_/D sky130_fd_sc_hd__o21a_1
XFILLER_164_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13090_ _13041_/S _12881_/X _13089_/X vssd1 vssd1 vccd1 vccd1 _13090_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12041_ _17798_/Q _12051_/B vssd1 vssd1 vccd1 vccd1 _12041_/X sky130_fd_sc_hd__or2_1
Xfanout1703 _08844_/Y vssd1 vssd1 vccd1 vccd1 _09457_/A sky130_fd_sc_hd__buf_12
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1714 _08828_/Y vssd1 vssd1 vccd1 vccd1 _12482_/S sky130_fd_sc_hd__buf_6
XFILLER_77_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1725 _08828_/A vssd1 vssd1 vccd1 vccd1 _16852_/A sky130_fd_sc_hd__buf_6
Xfanout1736 _18339_/Q vssd1 vssd1 vccd1 vccd1 _09657_/S sky130_fd_sc_hd__buf_12
XFILLER_104_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1747 _18117_/Q vssd1 vssd1 vccd1 vccd1 _14238_/A sky130_fd_sc_hd__buf_12
Xfanout760 _09160_/X vssd1 vssd1 vccd1 vccd1 _16470_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout1758 _09099_/A vssd1 vssd1 vccd1 vccd1 _09553_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout771 _17687_/S vssd1 vssd1 vccd1 vccd1 _17689_/S sky130_fd_sc_hd__clkbuf_16
X_15800_ _18593_/Q _15800_/A2 _15794_/Y _15799_/Y _17376_/A vssd1 vssd1 vccd1 vccd1
+ _18593_/D sky130_fd_sc_hd__o221a_1
Xfanout1769 _10471_/S vssd1 vssd1 vccd1 vccd1 _10866_/S sky130_fd_sc_hd__buf_4
Xfanout782 _16586_/S vssd1 vssd1 vccd1 vccd1 _16589_/S sky130_fd_sc_hd__buf_12
X_16780_ _19281_/Q _16783_/C _16780_/B1 vssd1 vssd1 vccd1 vccd1 _16780_/Y sky130_fd_sc_hd__o21ai_1
X_13992_ _17961_/Q _14028_/A vssd1 vssd1 vccd1 vccd1 _13992_/X sky130_fd_sc_hd__or2_1
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout793 _16352_/S vssd1 vssd1 vccd1 vccd1 _16358_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ _15729_/X _15730_/Y _15731_/B1 vssd1 vssd1 vccd1 vccd1 _15731_/Y sky130_fd_sc_hd__o21ai_1
X_12943_ _12794_/X _12797_/X _12943_/S vssd1 vssd1 vccd1 vccd1 _12943_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18450_ _18884_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _18587_/Q _18586_/Q _15662_/C vssd1 vssd1 vccd1 vccd1 _15704_/C sky130_fd_sc_hd__and3_2
X_12874_ _12678_/X _12726_/A _12942_/S vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__mux2_1
XANTENNA_120 _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _11814_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 _11853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17401_ _11732_/Y _15118_/A _15117_/A _17792_/Q _15116_/B vssd1 vssd1 vccd1 vccd1
+ _17401_/X sky130_fd_sc_hd__a221o_1
X_14613_ _17672_/A0 _18420_/Q _14630_/S vssd1 vssd1 vccd1 vccd1 _18420_/D sky130_fd_sc_hd__mux2_1
XANTENNA_153 _11872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11825_ _11846_/A _11825_/B vssd1 vssd1 vccd1 vccd1 _11826_/B sky130_fd_sc_hd__nor2_1
XFILLER_221_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_164 _13976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18381_ _19466_/CLK _18381_/D vssd1 vssd1 vccd1 vccd1 _18381_/Q sky130_fd_sc_hd__dfxtp_4
X_15593_ _15782_/A1 _15592_/X _15782_/B1 vssd1 vssd1 vccd1 vccd1 _15593_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _14000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 _13659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_197 _13886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17332_ _17342_/A _17332_/B vssd1 vssd1 vccd1 vccd1 _19463_/D sky130_fd_sc_hd__and2_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14596_/A _14544_/B vssd1 vssd1 vccd1 vccd1 _18380_/D sky130_fd_sc_hd__or2_1
XFILLER_230_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _18574_/Q _11759_/A2 _11844_/A _11683_/B vssd1 vssd1 vccd1 vccd1 _11756_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10707_ _10707_/A _10707_/B vssd1 vssd1 vccd1 vccd1 _10707_/X sky130_fd_sc_hd__or2_1
XFILLER_230_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14475_ _18327_/Q _17679_/A0 _14486_/S vssd1 vssd1 vccd1 vccd1 _18327_/D sky130_fd_sc_hd__mux2_1
X_17263_ _18115_/Q _17129_/A _17462_/A _17244_/B vssd1 vssd1 vccd1 vccd1 _17263_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11687_ _11687_/A _11774_/B vssd1 vssd1 vccd1 vccd1 _11687_/Y sky130_fd_sc_hd__nor2_2
XFILLER_186_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19002_ _19163_/CLK _19002_/D vssd1 vssd1 vccd1 vccd1 _19002_/Q sky130_fd_sc_hd__dfxtp_1
X_13426_ input270/X _12536_/Y _13847_/A2 _17870_/Q vssd1 vssd1 vccd1 vccd1 _13426_/X
+ sky130_fd_sc_hd__a22o_1
X_16214_ _17678_/A0 _18830_/Q _16226_/S vssd1 vssd1 vccd1 vccd1 _18830_/D sky130_fd_sc_hd__mux2_1
X_17194_ _19416_/Q fanout533/X _17513_/A _17119_/B vssd1 vssd1 vccd1 vccd1 _17195_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_10638_ _10532_/A _17682_/A0 _10637_/Y _11800_/B vssd1 vssd1 vccd1 vccd1 _11869_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16145_ _18775_/Q _16145_/B _16145_/C vssd1 vssd1 vccd1 vccd1 _16145_/X sky130_fd_sc_hd__or3_1
X_13357_ _14155_/B _12756_/Y _13357_/S vssd1 vssd1 vccd1 vccd1 _13357_/X sky130_fd_sc_hd__mux2_1
X_10569_ _10662_/A1 _19578_/Q _10645_/S _19610_/Q _10668_/S vssd1 vssd1 vccd1 vccd1
+ _10569_/X sky130_fd_sc_hd__o221a_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12308_ _14688_/A _12308_/B _16819_/A _16819_/B vssd1 vssd1 vccd1 vccd1 _12308_/X
+ sky130_fd_sc_hd__or4_1
X_16076_ _16074_/X _16075_/Y _16070_/Y vssd1 vssd1 vccd1 vccd1 _16076_/X sky130_fd_sc_hd__a21o_1
X_13288_ _13438_/A _13274_/Y _13563_/B1 vssd1 vssd1 vccd1 vccd1 _13289_/B sky130_fd_sc_hd__a21oi_1
X_15027_ _18516_/Q input193/X _15038_/S vssd1 vssd1 vccd1 vccd1 _18516_/D sky130_fd_sc_hd__mux2_1
X_12239_ _17878_/Q _12240_/C _17879_/Q vssd1 vssd1 vccd1 vccd1 _12241_/B sky130_fd_sc_hd__a21oi_1
XFILLER_269_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16978_ _16981_/B _17591_/C _16824_/A vssd1 vssd1 vccd1 vccd1 _17217_/B sky130_fd_sc_hd__or3b_4
XFILLER_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput4 coreIndex[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_6
X_18717_ _19142_/CLK _18717_/D vssd1 vssd1 vccd1 vccd1 _18717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15929_ input2/X input268/X _15947_/S vssd1 vssd1 vccd1 vccd1 _15929_/X sky130_fd_sc_hd__mux2_1
XFILLER_265_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09450_ _10263_/A1 _17765_/Q _09464_/S _18314_/Q _10264_/S vssd1 vssd1 vccd1 vccd1
+ _09450_/X sky130_fd_sc_hd__o221a_1
XFILLER_64_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18648_ _19211_/CLK _18648_/D vssd1 vssd1 vccd1 vccd1 _18648_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09381_ _09379_/X _09380_/X _09381_/S vssd1 vssd1 vccd1 vccd1 _09381_/X sky130_fd_sc_hd__mux2_1
XFILLER_212_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18579_ _19507_/CLK _18579_/D vssd1 vssd1 vccd1 vccd1 _18579_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput330 _11747_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[7] sky130_fd_sc_hd__buf_4
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput341 _11840_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[16] sky130_fd_sc_hd__buf_4
Xoutput352 _11886_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[26] sky130_fd_sc_hd__buf_4
XFILLER_273_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput363 _11802_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[7] sky130_fd_sc_hd__buf_4
Xoutput374 _11705_/Y vssd1 vssd1 vccd1 vccd1 csb1[0] sky130_fd_sc_hd__buf_4
XFILLER_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput385 _11938_/X vssd1 vssd1 vccd1 vccd1 din0[18] sky130_fd_sc_hd__buf_4
XFILLER_160_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput396 _11948_/X vssd1 vssd1 vccd1 vccd1 din0[28] sky130_fd_sc_hd__buf_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09717_ _18536_/Q _18411_/Q _10717_/S vssd1 vssd1 vccd1 vccd1 _09717_/X sky130_fd_sc_hd__mux2_1
XFILLER_216_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09648_ _13044_/S _09648_/B vssd1 vssd1 vccd1 vccd1 _13033_/A sky130_fd_sc_hd__or2_1
XFILLER_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09579_ _10742_/A1 _09578_/X _09577_/X vssd1 vssd1 vccd1 vccd1 _09579_/X sky130_fd_sc_hd__o21a_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11610_ _18563_/Q _18438_/Q _11613_/S vssd1 vssd1 vccd1 vccd1 _11610_/X sky130_fd_sc_hd__mux2_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12590_ _12453_/X _13930_/A1 _13253_/B1 vssd1 vssd1 vccd1 vccd1 _12590_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_212_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11541_ _11541_/A _11541_/B vssd1 vssd1 vccd1 vccd1 _13697_/A sky130_fd_sc_hd__nor2_8
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14260_ _18128_/Q _14260_/B vssd1 vssd1 vccd1 vccd1 _14260_/X sky130_fd_sc_hd__or2_1
XFILLER_128_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11472_ _11481_/A _19175_/Q _11472_/C vssd1 vssd1 vccd1 vccd1 _11472_/X sky130_fd_sc_hd__and3_1
XFILLER_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13211_ _19433_/Q _12560_/B _13209_/X _13210_/X _12560_/A vssd1 vssd1 vccd1 vccd1
+ _13211_/X sky130_fd_sc_hd__o221a_1
X_10423_ _18074_/Q _10364_/B _10422_/X _10419_/S vssd1 vssd1 vccd1 vccd1 _10423_/X
+ sky130_fd_sc_hd__o211a_1
X_14191_ _16964_/A _14191_/B vssd1 vssd1 vccd1 vccd1 _18093_/D sky130_fd_sc_hd__and2_1
XFILLER_164_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13142_ _13896_/B2 _13137_/Y _13140_/X _12732_/S _13141_/Y vssd1 vssd1 vccd1 vccd1
+ _13142_/X sky130_fd_sc_hd__o221a_4
XFILLER_100_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10354_ _10354_/A1 _18231_/Q _10353_/S _18966_/Q _10205_/S vssd1 vssd1 vccd1 vccd1
+ _10354_/X sky130_fd_sc_hd__o221a_1
XFILLER_151_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13073_ _17861_/Q _13945_/A2 _13061_/X _13303_/B2 _13952_/B1 vssd1 vssd1 vccd1 vccd1
+ _13073_/X sky130_fd_sc_hd__a221o_1
X_17950_ _18627_/CLK _17950_/D vssd1 vssd1 vccd1 vccd1 _17950_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10285_ _11199_/S1 _10275_/X _10284_/X _11516_/B1 vssd1 vssd1 vccd1 vccd1 _10285_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16901_ _18756_/Q _16961_/A2 _16969_/B1 input220/X _16969_/C1 vssd1 vssd1 vccd1 vccd1
+ _16901_/X sky130_fd_sc_hd__a221o_1
XFILLER_151_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1500 _09498_/S vssd1 vssd1 vccd1 vccd1 _09883_/B sky130_fd_sc_hd__buf_6
X_12024_ _12024_/A _17724_/B vssd1 vssd1 vccd1 vccd1 _12024_/Y sky130_fd_sc_hd__nand2_2
Xfanout1511 _10199_/S vssd1 vssd1 vccd1 vccd1 _10353_/S sky130_fd_sc_hd__buf_6
XFILLER_250_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1522 _10426_/S vssd1 vssd1 vccd1 vccd1 _11503_/S0 sky130_fd_sc_hd__buf_6
X_17881_ _19323_/CLK _17881_/D vssd1 vssd1 vccd1 vccd1 _17881_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1533 _10275_/S vssd1 vssd1 vccd1 vccd1 _09718_/S sky130_fd_sc_hd__buf_6
XFILLER_39_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1544 _10649_/A1 vssd1 vssd1 vccd1 vccd1 _10668_/S sky130_fd_sc_hd__buf_8
X_19620_ _19620_/CLK _19620_/D vssd1 vssd1 vccd1 vccd1 _19620_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1555 _09381_/S vssd1 vssd1 vccd1 vccd1 _10225_/S sky130_fd_sc_hd__buf_6
X_16832_ _16821_/A _17815_/Q _12486_/X vssd1 vssd1 vccd1 vccd1 _17051_/B sky130_fd_sc_hd__a21o_1
Xfanout1566 _11279_/B1 vssd1 vssd1 vccd1 vccd1 _11623_/A1 sky130_fd_sc_hd__buf_6
XFILLER_266_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1577 fanout1581/X vssd1 vssd1 vccd1 vccd1 _08967_/S sky130_fd_sc_hd__buf_4
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1588 _10211_/A1 vssd1 vssd1 vccd1 vccd1 _09978_/A1 sky130_fd_sc_hd__buf_8
Xfanout590 _12073_/B vssd1 vssd1 vccd1 vccd1 _12087_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_281_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1599 _11516_/B1 vssd1 vssd1 vccd1 vccd1 _11438_/B1 sky130_fd_sc_hd__buf_8
XFILLER_219_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19551_ _19553_/CLK _19551_/D vssd1 vssd1 vccd1 vccd1 _19551_/Q sky130_fd_sc_hd__dfxtp_1
X_16763_ _16768_/A _16763_/B _16767_/C vssd1 vssd1 vccd1 vccd1 _19274_/D sky130_fd_sc_hd__nor3_1
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13975_ _14033_/A1 _12550_/X _13974_/X _14037_/C1 vssd1 vssd1 vccd1 vccd1 _17952_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18502_ _19286_/CLK _18502_/D vssd1 vssd1 vccd1 vccd1 _18502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15714_ _15696_/A _15693_/Y _15695_/B vssd1 vssd1 vccd1 vccd1 _15715_/B sky130_fd_sc_hd__o21ai_2
XFILLER_262_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19482_ _19482_/CLK _19482_/D vssd1 vssd1 vccd1 vccd1 _19482_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ _14714_/A _12868_/B _18104_/Q vssd1 vssd1 vccd1 vccd1 _12927_/B sky130_fd_sc_hd__o21ba_1
X_16694_ _19250_/Q _16699_/D _19251_/Q vssd1 vssd1 vccd1 vccd1 _16696_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18433_ _19565_/CLK _18433_/D vssd1 vssd1 vccd1 vccd1 _18433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_261_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15645_ _15645_/A _15645_/B vssd1 vssd1 vccd1 vccd1 _15645_/X sky130_fd_sc_hd__or2_2
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12857_ _19488_/Q _12856_/X _12857_/S vssd1 vssd1 vccd1 vccd1 _12857_/X sky130_fd_sc_hd__mux2_2
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18364_ _19642_/CLK _18364_/D vssd1 vssd1 vccd1 vccd1 _18364_/Q sky130_fd_sc_hd__dfxtp_1
X_11808_ _11808_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__or2_4
X_15576_ _15787_/A _15639_/A vssd1 vssd1 vccd1 vccd1 _15576_/X sky130_fd_sc_hd__or2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _18102_/Q _12788_/B vssd1 vssd1 vccd1 vccd1 _12789_/B sky130_fd_sc_hd__and2_1
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17313_/Y _17314_/X _16048_/A vssd1 vssd1 vccd1 vccd1 _19455_/D sky130_fd_sc_hd__a21oi_1
XFILLER_202_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14527_ _18405_/Q _14527_/B vssd1 vssd1 vccd1 vccd1 _14527_/Y sky130_fd_sc_hd__nor2_1
X_11739_ _11739_/A _11739_/B vssd1 vssd1 vccd1 vccd1 _11740_/A sky130_fd_sc_hd__xnor2_4
X_18295_ _18593_/CLK _18295_/D vssd1 vssd1 vccd1 vccd1 _18295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17246_ _17244_/Y _17245_/X _17255_/A vssd1 vssd1 vccd1 vccd1 _19432_/D sky130_fd_sc_hd__a21oi_1
X_14458_ _18310_/Q _16595_/A0 _14486_/S vssd1 vssd1 vccd1 vccd1 _18310_/D sky130_fd_sc_hd__mux2_1
X_13409_ _13443_/B _13961_/A vssd1 vssd1 vccd1 vccd1 _13409_/Y sky130_fd_sc_hd__nand2_1
X_14389_ _16431_/A1 _18240_/Q _14412_/S vssd1 vssd1 vccd1 vccd1 _18240_/D sky130_fd_sc_hd__mux2_1
X_17177_ _17285_/A _17177_/B vssd1 vssd1 vccd1 vccd1 _19410_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16128_ _16140_/A1 _16127_/Y _16128_/B1 vssd1 vssd1 vccd1 vccd1 _18766_/D sky130_fd_sc_hd__a21oi_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08950_ _08950_/A _16392_/C vssd1 vssd1 vccd1 vccd1 _08950_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_170_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16059_ _08861_/Y _16053_/Y _16056_/Y _16058_/X vssd1 vssd1 vccd1 vccd1 _16059_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08881_ _09854_/A _08882_/B vssd1 vssd1 vccd1 vccd1 _08881_/X sky130_fd_sc_hd__and2_4
XFILLER_285_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09502_ _18445_/Q _18346_/Q _09883_/B vssd1 vssd1 vccd1 vccd1 _09502_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09433_ _17959_/Q _11216_/A2 _09017_/X _11687_/A vssd1 vssd1 vccd1 vccd1 _09433_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09364_ _11452_/A _09334_/X _09363_/X vssd1 vssd1 vccd1 vccd1 _11804_/A sky130_fd_sc_hd__o21ai_4
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_20 _14960_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ _09293_/X _09294_/X _09374_/S vssd1 vssd1 vccd1 vccd1 _09295_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 _17214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_42 _12600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 _09743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_64 _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_86 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_97 _13515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__nand2_2
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ _13294_/A _13761_/A _13968_/A1 _13759_/X vssd1 vssd1 vccd1 vccd1 _13760_/X
+ sky130_fd_sc_hd__o211a_1
X_10972_ _11360_/A1 _18326_/Q _17777_/Q _11340_/B2 vssd1 vssd1 vccd1 vccd1 _10972_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12711_ _12614_/B _12648_/B _12732_/S vssd1 vssd1 vccd1 vccd1 _12711_/X sky130_fd_sc_hd__mux2_1
XFILLER_271_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13691_ _13747_/B2 _13680_/X _13690_/X vssd1 vssd1 vccd1 vccd1 _13691_/X sky130_fd_sc_hd__a21o_4
XFILLER_188_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12642_ _13616_/A _13615_/B _12640_/Y vssd1 vssd1 vccd1 vccd1 _12643_/B sky130_fd_sc_hd__o21ai_1
X_15430_ _15432_/A _15432_/B vssd1 vssd1 vccd1 vccd1 _15430_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15361_ _15361_/A _15361_/B vssd1 vssd1 vccd1 vccd1 _15456_/A sky130_fd_sc_hd__xor2_2
X_12573_ _12577_/A _12584_/B vssd1 vssd1 vccd1 vccd1 _12576_/B sky130_fd_sc_hd__or2_2
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17100_ _17190_/B _17116_/A2 _17099_/X _17106_/C1 vssd1 vssd1 vccd1 vccd1 _19383_/D
+ sky130_fd_sc_hd__o211a_1
X_14312_ _18169_/Q _16431_/A1 _14335_/S vssd1 vssd1 vccd1 vccd1 _18169_/D sky130_fd_sc_hd__mux2_1
X_11524_ _13311_/A vssd1 vssd1 vccd1 vccd1 _11681_/A sky130_fd_sc_hd__clkinv_4
X_18080_ _19650_/CLK _18080_/D vssd1 vssd1 vccd1 vccd1 _18080_/Q sky130_fd_sc_hd__dfxtp_1
X_15292_ _18571_/Q _15314_/C vssd1 vssd1 vccd1 vccd1 _15292_/X sky130_fd_sc_hd__xor2_1
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14243_ _18293_/Q _14267_/A2 _14242_/X _14452_/B vssd1 vssd1 vccd1 vccd1 _18119_/D
+ sky130_fd_sc_hd__o211a_1
X_17031_ _19352_/Q _17041_/B vssd1 vssd1 vccd1 vccd1 _17031_/X sky130_fd_sc_hd__or2_1
X_11455_ _18638_/Q _18060_/Q _11455_/S vssd1 vssd1 vccd1 vccd1 _11455_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10406_ _11458_/A1 _18230_/Q _11379_/S _18965_/Q vssd1 vssd1 vccd1 vccd1 _10406_/X
+ sky130_fd_sc_hd__o22a_1
X_14174_ _18698_/Q _18085_/Q _14186_/S vssd1 vssd1 vccd1 vccd1 _14175_/B sky130_fd_sc_hd__mux2_1
XFILLER_171_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11386_ _18029_/Q _17997_/Q _11386_/S vssd1 vssd1 vccd1 vccd1 _11386_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13125_ _13125_/A _13349_/B vssd1 vssd1 vccd1 vccd1 _13125_/X sky130_fd_sc_hd__and2_1
X_10337_ _18653_/Q _18075_/Q _19094_/Q _18998_/Q _09179_/B _10337_/S1 vssd1 vssd1
+ vccd1 vccd1 _10337_/X sky130_fd_sc_hd__mux4_1
X_18982_ _19076_/CLK _18982_/D vssd1 vssd1 vccd1 vccd1 _18982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17933_ _18749_/CLK _17933_/D vssd1 vssd1 vccd1 vccd1 _17933_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13159_/C _13056_/B vssd1 vssd1 vccd1 vccd1 _13056_/X sky130_fd_sc_hd__or2_2
X_10268_ _10265_/X _10267_/X _10180_/A vssd1 vssd1 vccd1 vccd1 _10268_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1330 _10707_/A vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__buf_6
XFILLER_94_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12007_ _17774_/Q _17708_/A0 _12013_/S vssd1 vssd1 vccd1 vccd1 _17774_/D sky130_fd_sc_hd__mux2_1
XFILLER_267_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1341 _10618_/S vssd1 vssd1 vccd1 vccd1 _11577_/S sky130_fd_sc_hd__buf_8
XFILLER_266_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1352 _09914_/C1 vssd1 vssd1 vccd1 vccd1 _11478_/S sky130_fd_sc_hd__buf_6
X_17864_ _17865_/CLK _17864_/D vssd1 vssd1 vccd1 vccd1 _17864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10199_ _18561_/Q _18436_/Q _10199_/S vssd1 vssd1 vccd1 vccd1 _10199_/X sky130_fd_sc_hd__mux2_1
XFILLER_266_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1363 _10864_/S vssd1 vssd1 vccd1 vccd1 _11576_/S sky130_fd_sc_hd__buf_6
XFILLER_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_159_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19537_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_239_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1374 _09843_/S vssd1 vssd1 vccd1 vccd1 _10467_/S sky130_fd_sc_hd__buf_4
X_19603_ _19635_/CLK _19603_/D vssd1 vssd1 vccd1 vccd1 _19603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16815_ _19294_/Q _19293_/Q _16815_/C vssd1 vssd1 vccd1 vccd1 _16816_/C sky130_fd_sc_hd__nand3_2
Xfanout1385 fanout1386/X vssd1 vssd1 vccd1 vccd1 _11154_/S sky130_fd_sc_hd__buf_4
Xfanout1396 _10249_/S vssd1 vssd1 vccd1 vccd1 _09464_/S sky130_fd_sc_hd__buf_6
XFILLER_266_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17795_ _19650_/CLK _17795_/D vssd1 vssd1 vccd1 vccd1 _17795_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19534_ _19534_/CLK _19534_/D vssd1 vssd1 vccd1 vccd1 _19534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16746_ _19268_/Q _16746_/B vssd1 vssd1 vccd1 vccd1 _16751_/C sky130_fd_sc_hd__and2_2
XFILLER_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13958_ _13958_/A _13958_/B vssd1 vssd1 vccd1 vccd1 _13958_/X sky130_fd_sc_hd__or2_1
XFILLER_81_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12909_ input283/X _12851_/B _12859_/S vssd1 vssd1 vccd1 vccd1 _12909_/X sky130_fd_sc_hd__a21o_1
XFILLER_262_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19465_ _19465_/CLK _19465_/D vssd1 vssd1 vccd1 vccd1 _19465_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_262_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16677_ _16677_/A _16677_/B _16677_/C _16677_/D vssd1 vssd1 vccd1 vccd1 _16688_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13889_ _13289_/A _13887_/Y _13888_/X _13904_/B _13294_/A vssd1 vssd1 vccd1 vccd1
+ _13889_/X sky130_fd_sc_hd__o32a_1
X_18416_ _19595_/CLK _18416_/D vssd1 vssd1 vccd1 vccd1 _18416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15628_ _19479_/Q _19413_/Q vssd1 vssd1 vccd1 vccd1 _15628_/X sky130_fd_sc_hd__and2_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19396_ _19526_/CLK _19396_/D vssd1 vssd1 vccd1 vccd1 _19396_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_222_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18347_ _19625_/CLK _18347_/D vssd1 vssd1 vccd1 vccd1 _18347_/Q sky130_fd_sc_hd__dfxtp_1
X_15559_ _15556_/X _15558_/X _15638_/A vssd1 vssd1 vccd1 vccd1 _15580_/B sky130_fd_sc_hd__a21oi_4
XFILLER_175_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09080_ _12443_/A _09080_/B _09080_/C vssd1 vssd1 vccd1 vccd1 _13916_/A sky130_fd_sc_hd__or3_4
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18278_ _18734_/CLK _18278_/D vssd1 vssd1 vccd1 vccd1 _18278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput40 core_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_2
X_17229_ _18104_/Q _17219_/A _17129_/Y _17219_/B vssd1 vssd1 vccd1 vccd1 _17229_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 dout0[17] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput62 dout0[27] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_2
Xinput73 dout0[37] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_2
Xinput84 dout0[47] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_2
Xinput95 dout0[57] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09982_ _09984_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _12838_/S sky130_fd_sc_hd__and2b_2
XFILLER_116_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08933_ _12053_/A _08995_/B _08932_/X _17820_/Q vssd1 vssd1 vccd1 vccd1 _08933_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_254_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08864_ _18080_/Q _17887_/Q vssd1 vssd1 vccd1 vccd1 _08864_/X sky130_fd_sc_hd__and2b_1
XFILLER_112_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09416_ _10275_/S _09415_/X _08903_/A vssd1 vssd1 vccd1 vccd1 _09416_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09347_ _09340_/X _09346_/X _09337_/X _09343_/X _08843_/A _12408_/A vssd1 vssd1 vccd1
+ vccd1 _09347_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ _11452_/A _16204_/A0 _09277_/X vssd1 vssd1 vccd1 vccd1 _11808_/A sky130_fd_sc_hd__o21ai_4
XFILLER_166_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ _11238_/X _11239_/X _11248_/S vssd1 vssd1 vccd1 vccd1 _11240_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11171_ _18859_/Q _18891_/Q _11171_/S vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10122_ _12442_/A _11490_/B _11489_/B1 _10121_/Y vssd1 vssd1 vccd1 vccd1 _10159_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14930_ _18494_/Q _15011_/A2 _14929_/Y _16787_/A vssd1 vssd1 vccd1 vccd1 _18494_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_88_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10053_ _10033_/S _10052_/X _10051_/X _11274_/S1 vssd1 vssd1 vccd1 vccd1 _10053_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14861_ _17807_/Q _15002_/B vssd1 vssd1 vccd1 vccd1 _14861_/X sky130_fd_sc_hd__or2_1
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16600_ _17700_/A0 _19203_/Q _16622_/S vssd1 vssd1 vccd1 vccd1 _19203_/D sky130_fd_sc_hd__mux2_1
XFILLER_264_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _13812_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _14152_/A sky130_fd_sc_hd__xnor2_4
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17580_ _19532_/Q _17561_/B _17588_/B1 _17579_/X vssd1 vssd1 vccd1 vccd1 _19532_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14792_ _18111_/Q _14994_/B _14771_/X _14791_/X vssd1 vssd1 vccd1 vccd1 _14792_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16531_ _17664_/A0 _19136_/Q _16548_/S vssd1 vssd1 vccd1 vccd1 _19136_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13743_ _13743_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13758_/B sky130_fd_sc_hd__or2_1
X_10955_ _10953_/X _10954_/X _11361_/S vssd1 vssd1 vccd1 vccd1 _10955_/X sky130_fd_sc_hd__mux2_1
XFILLER_244_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19250_ _19295_/CLK _19250_/D vssd1 vssd1 vccd1 vccd1 _19250_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16462_ _16462_/A0 _19069_/Q _16485_/S vssd1 vssd1 vccd1 vccd1 _19069_/D sky130_fd_sc_hd__mux2_1
X_13674_ _15133_/A _13672_/X _13673_/Y _13869_/B2 vssd1 vssd1 vccd1 vccd1 _13675_/B
+ sky130_fd_sc_hd__a22o_1
X_10886_ _10040_/S _10885_/X _11623_/A1 vssd1 vssd1 vccd1 vccd1 _10887_/B sky130_fd_sc_hd__a21o_1
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18201_ _18201_/CLK _18201_/D vssd1 vssd1 vccd1 vccd1 _18201_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15413_ _18576_/Q _15412_/B _15437_/B1 vssd1 vssd1 vccd1 vccd1 _15414_/B sky130_fd_sc_hd__o21ai_1
X_19181_ _19213_/CLK _19181_/D vssd1 vssd1 vccd1 vccd1 _19181_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12625_ _12625_/A _12625_/B vssd1 vssd1 vccd1 vccd1 _12625_/Y sky130_fd_sc_hd__nor2_1
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16393_ _16393_/A _16591_/B vssd1 vssd1 vccd1 vccd1 _16393_/Y sky130_fd_sc_hd__nand2_2
XFILLER_31_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18132_ _19444_/CLK _18132_/D vssd1 vssd1 vccd1 vccd1 _18132_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12556_ _12768_/B _12561_/B vssd1 vssd1 vccd1 vccd1 _12556_/Y sky130_fd_sc_hd__nor2_1
X_15344_ _19435_/Q _15411_/B _17211_/A _15343_/Y vssd1 vssd1 vccd1 vccd1 _15344_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ _11505_/X _11506_/X _11507_/S vssd1 vssd1 vccd1 vccd1 _11507_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18063_ _19586_/CLK _18063_/D vssd1 vssd1 vccd1 vccd1 _18063_/Q sky130_fd_sc_hd__dfxtp_1
X_12487_ _12488_/A _17913_/Q _12486_/X vssd1 vssd1 vccd1 vccd1 _12572_/B sky130_fd_sc_hd__a21o_1
X_15275_ _19464_/Q _19398_/Q vssd1 vssd1 vccd1 vccd1 _15275_/Y sky130_fd_sc_hd__nor2_2
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17014_ _17589_/A _17032_/A2 _17013_/X _17360_/A vssd1 vssd1 vccd1 vccd1 _19343_/D
+ sky130_fd_sc_hd__o211a_1
X_11438_ _11433_/Y _11437_/Y _11438_/B1 vssd1 vssd1 vccd1 vccd1 _11438_/X sky130_fd_sc_hd__a21o_1
X_14226_ _18111_/Q _14244_/B vssd1 vssd1 vccd1 vccd1 _14226_/X sky130_fd_sc_hd__or2_1
XFILLER_256_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14157_ _12440_/X _14155_/A _14155_/Y _14156_/X vssd1 vssd1 vccd1 vccd1 _14158_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_259_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11369_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _12626_/B sky130_fd_sc_hd__nor2_4
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13108_ _19497_/Q _13064_/B _13243_/B1 _13107_/X vssd1 vssd1 vccd1 vccd1 _13108_/X
+ sky130_fd_sc_hd__o211a_1
X_18965_ _19157_/CLK _18965_/D vssd1 vssd1 vccd1 vccd1 _18965_/Q sky130_fd_sc_hd__dfxtp_1
X_14088_ _17671_/A0 _18028_/Q _14106_/S vssd1 vssd1 vccd1 vccd1 _18028_/D sky130_fd_sc_hd__mux2_1
XFILLER_224_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17916_ _18881_/CLK _17916_/D vssd1 vssd1 vccd1 vccd1 _17916_/Q sky130_fd_sc_hd__dfxtp_4
X_13039_ _12795_/X _12806_/X _13039_/S vssd1 vssd1 vccd1 vccd1 _13039_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18896_ _19607_/CLK _18896_/D vssd1 vssd1 vccd1 vccd1 _18896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1160 _16005_/A2 vssd1 vssd1 vccd1 vccd1 _16019_/A2 sky130_fd_sc_hd__buf_4
XFILLER_39_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1171 _15946_/A2 vssd1 vssd1 vccd1 vccd1 _15949_/A2 sky130_fd_sc_hd__buf_4
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17847_ _19324_/CLK _17847_/D vssd1 vssd1 vccd1 vccd1 _17847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1182 _15404_/B vssd1 vssd1 vccd1 vccd1 _15304_/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1193 _15953_/Y vssd1 vssd1 vccd1 vccd1 _16002_/B1 sky130_fd_sc_hd__buf_4
XFILLER_226_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17778_ _19649_/CLK _17778_/D vssd1 vssd1 vccd1 vccd1 _17778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19517_ _19546_/CLK _19517_/D vssd1 vssd1 vccd1 vccd1 _19517_/Q sky130_fd_sc_hd__dfxtp_1
X_16729_ _19262_/Q _19261_/Q _16729_/C vssd1 vssd1 vccd1 vccd1 _16736_/D sky130_fd_sc_hd__and3_1
XFILLER_223_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19448_ _19448_/CLK _19448_/D vssd1 vssd1 vccd1 vccd1 _19448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09201_ _09197_/X _09198_/X _10225_/S vssd1 vssd1 vccd1 vccd1 _09201_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19379_ _19542_/CLK _19379_/D vssd1 vssd1 vccd1 vccd1 _19379_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_56_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19648_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_188_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09132_ _19110_/Q _19142_/Q _11455_/S vssd1 vssd1 vccd1 vccd1 _09132_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09063_ _17900_/Q _12264_/A vssd1 vssd1 vccd1 vccd1 _12754_/B sky130_fd_sc_hd__nor2_2
XFILLER_190_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09965_ _18308_/Q _17759_/Q _09966_/S vssd1 vssd1 vccd1 vccd1 _09965_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08916_ _12089_/A _17801_/Q vssd1 vssd1 vccd1 vccd1 _16392_/C sky130_fd_sc_hd__and2_4
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _12602_/B vssd1 vssd1 vccd1 vccd1 _09896_/Y sky130_fd_sc_hd__inv_2
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _17906_/Q vssd1 vssd1 vccd1 vccd1 _08897_/A sky130_fd_sc_hd__inv_2
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_505 _08874_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_516 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_527 _11132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_538 input233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_549 _12320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10740_ _10737_/X _10738_/X _10739_/X _10742_/A1 _10746_/S vssd1 vssd1 vccd1 vccd1
+ _10740_/X sky130_fd_sc_hd__a221o_1
XFILLER_159_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10671_ _11602_/C1 _10664_/X _11286_/B1 vssd1 vssd1 vccd1 vccd1 _10671_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_167_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _17887_/Q _12433_/B _12409_/X _12408_/X _13981_/C1 vssd1 vssd1 vccd1 vccd1
+ _17911_/D sky130_fd_sc_hd__o311a_1
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13390_ _12833_/Y _13389_/X _13390_/S vssd1 vssd1 vccd1 vccd1 _13390_/X sky130_fd_sc_hd__mux2_1
XFILLER_223_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12341_ _17888_/Q _12382_/A _12340_/Y _12383_/C1 vssd1 vssd1 vccd1 vccd1 _17888_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_166_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15060_ _18544_/Q _17671_/A0 _15076_/S vssd1 vssd1 vccd1 vccd1 _18544_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ _18775_/Q _16143_/C _18776_/Q vssd1 vssd1 vccd1 vccd1 _12272_/X sky130_fd_sc_hd__and3b_2
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14011_ _14033_/A1 _13527_/X _14010_/X _14029_/C1 vssd1 vssd1 vccd1 vccd1 _17970_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11223_ _17935_/Q _08948_/B _11222_/X _08947_/B vssd1 vssd1 vccd1 vccd1 _11223_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11154_ _18032_/Q _18000_/Q _11154_/S vssd1 vssd1 vccd1 vccd1 _11154_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10105_ _10243_/A _10100_/X _10102_/X _10104_/X _09264_/S vssd1 vssd1 vccd1 vccd1
+ _10105_/Y sky130_fd_sc_hd__o221ai_4
X_18750_ _18775_/CLK _18750_/D vssd1 vssd1 vccd1 vccd1 _18750_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15962_ _18696_/Q _15970_/A2 _15976_/B1 _18745_/Q _15976_/C1 vssd1 vssd1 vccd1 vccd1
+ _15962_/X sky130_fd_sc_hd__a221o_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11085_ _19052_/Q _19020_/Q _11094_/S vssd1 vssd1 vccd1 vccd1 _11085_/X sky130_fd_sc_hd__mux2_1
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput230 localMemory_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 input230/X sky130_fd_sc_hd__buf_12
XFILLER_283_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17701_ _17701_/A0 _19627_/Q _17719_/S vssd1 vssd1 vccd1 vccd1 _19627_/D sky130_fd_sc_hd__mux2_1
XFILLER_209_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput241 localMemory_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input241/X sky130_fd_sc_hd__buf_8
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput252 localMemory_wb_we_i vssd1 vssd1 vccd1 vccd1 input252/X sky130_fd_sc_hd__clkbuf_2
X_14913_ _14911_/X _14912_/X _14913_/B1 vssd1 vssd1 vccd1 vccd1 _14913_/X sky130_fd_sc_hd__a21o_1
X_10036_ _10034_/X _10035_/X _10036_/S vssd1 vssd1 vccd1 vccd1 _10036_/X sky130_fd_sc_hd__mux2_1
Xinput263 manufacturerID[9] vssd1 vssd1 vccd1 vccd1 _15884_/A sky130_fd_sc_hd__buf_4
X_18681_ _18683_/CLK _18681_/D vssd1 vssd1 vccd1 vccd1 _18681_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput274 partID[4] vssd1 vssd1 vccd1 vccd1 _15902_/A sky130_fd_sc_hd__clkbuf_2
X_15893_ _15893_/A _15905_/B _15905_/C vssd1 vssd1 vccd1 vccd1 _15893_/X sky130_fd_sc_hd__and3_1
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _17665_/A0 _19560_/Q _17654_/S vssd1 vssd1 vccd1 vccd1 _19560_/D sky130_fd_sc_hd__mux2_1
XFILLER_252_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ input49/X input84/X _14844_/S vssd1 vssd1 vccd1 vccd1 _14845_/A sky130_fd_sc_hd__mux2_2
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17563_ _17563_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17563_/X sky130_fd_sc_hd__or2_1
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14775_ _14775_/A vssd1 vssd1 vccd1 vccd1 _14775_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ _14074_/C _14272_/B vssd1 vssd1 vccd1 vccd1 _17625_/A sky130_fd_sc_hd__nor2_8
X_19302_ _19363_/CLK _19302_/D vssd1 vssd1 vccd1 vccd1 _19302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16514_ _16547_/A0 _19120_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _19120_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13726_ _13931_/A _13724_/Y _13725_/X _13740_/B _13294_/A vssd1 vssd1 vccd1 vccd1
+ _13726_/X sky130_fd_sc_hd__o32a_1
XFILLER_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17494_ _19510_/Q _17493_/B _17492_/X _17493_/Y _17356_/A vssd1 vssd1 vccd1 vccd1
+ _19510_/D sky130_fd_sc_hd__o221a_1
X_10938_ _11305_/A1 _18613_/Q _18184_/Q _10929_/S vssd1 vssd1 vccd1 vccd1 _10938_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19233_ _19268_/CLK _19233_/D vssd1 vssd1 vccd1 vccd1 _19233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16445_ _19053_/Q _16610_/A0 _16457_/S vssd1 vssd1 vccd1 vccd1 _19053_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10869_ _10848_/X _10851_/X _10868_/X vssd1 vssd1 vccd1 vccd1 _10869_/X sky130_fd_sc_hd__a21o_1
X_13657_ _19382_/Q _13951_/A2 _13655_/X _13656_/X _13951_/C1 vssd1 vssd1 vccd1 vccd1
+ _13657_/X sky130_fd_sc_hd__o221a_4
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19164_ _19626_/CLK _19164_/D vssd1 vssd1 vccd1 vccd1 _19164_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _12999_/S _09736_/B _12985_/B vssd1 vssd1 vccd1 vccd1 _12610_/A sky130_fd_sc_hd__a21o_1
XFILLER_158_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _16476_/A0 _18987_/Q _16385_/S vssd1 vssd1 vccd1 vccd1 _18987_/D sky130_fd_sc_hd__mux2_1
X_13588_ _19412_/Q _13948_/A2 _13948_/B1 vssd1 vssd1 vccd1 vccd1 _13588_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18115_ _19450_/CLK _18115_/D vssd1 vssd1 vccd1 vccd1 _18115_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_145_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15327_ _18572_/Q _15351_/A2 _15318_/Y _15326_/X _17469_/C1 vssd1 vssd1 vccd1 vccd1
+ _18572_/D sky130_fd_sc_hd__o221a_1
X_12539_ _15890_/A _12536_/Y _12538_/Y input280/X _12505_/Y vssd1 vssd1 vccd1 vccd1
+ _12539_/X sky130_fd_sc_hd__a221o_1
X_19095_ _19159_/CLK _19095_/D vssd1 vssd1 vccd1 vccd1 _19095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18046_ _19648_/CLK _18046_/D vssd1 vssd1 vccd1 vccd1 _18046_/Q sky130_fd_sc_hd__dfxtp_1
X_15258_ _17916_/Q _15369_/A vssd1 vssd1 vccd1 vccd1 _15262_/A sky130_fd_sc_hd__nand2_2
XFILLER_172_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14209_ _18276_/Q _14267_/A2 _14208_/X _14452_/B vssd1 vssd1 vccd1 vccd1 _18102_/D
+ sky130_fd_sc_hd__o211a_1
X_15189_ _15189_/A _15189_/B vssd1 vssd1 vccd1 vccd1 _15189_/Y sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_174_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19519_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_103_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18683_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09750_ _09746_/X _09749_/X _09750_/S vssd1 vssd1 vccd1 vccd1 _09750_/X sky130_fd_sc_hd__mux2_1
X_18948_ _19140_/CLK _18948_/D vssd1 vssd1 vccd1 vccd1 _18948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09681_ _10323_/A1 _19135_/Q _09925_/S _19103_/Q vssd1 vssd1 vccd1 vccd1 _09681_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18879_ _19138_/CLK _18879_/D vssd1 vssd1 vccd1 vccd1 _18879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09115_ _11465_/A1 _17769_/Q _11455_/S _18318_/Q _09135_/S vssd1 vssd1 vccd1 vccd1
+ _09115_/X sky130_fd_sc_hd__o221a_1
XFILLER_210_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09046_ _18202_/Q _09046_/B vssd1 vssd1 vccd1 vccd1 _09046_/Y sky130_fd_sc_hd__nand2_1
XFILLER_276_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1907 _14928_/B1 vssd1 vssd1 vccd1 vccd1 _14918_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout920 _16245_/S vssd1 vssd1 vccd1 vccd1 _16259_/S sky130_fd_sc_hd__buf_12
XFILLER_131_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout931 _15083_/Y vssd1 vssd1 vccd1 vccd1 _15117_/A sky130_fd_sc_hd__buf_6
XFILLER_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout942 _14994_/B vssd1 vssd1 vccd1 vccd1 _14801_/B sky130_fd_sc_hd__buf_4
XFILLER_38_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09948_ _18102_/Q _09948_/B vssd1 vssd1 vccd1 vccd1 _09948_/X sky130_fd_sc_hd__or2_1
Xfanout953 _14599_/X vssd1 vssd1 vccd1 vccd1 _14631_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout964 _14108_/Y vssd1 vssd1 vccd1 vccd1 _14137_/S sky130_fd_sc_hd__buf_8
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout975 _13527_/B1 vssd1 vssd1 vccd1 vccd1 _13928_/A1 sky130_fd_sc_hd__clkbuf_16
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout986 _13973_/A2 vssd1 vssd1 vccd1 vccd1 _13742_/A2 sky130_fd_sc_hd__clkbuf_8
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout997 _10459_/X vssd1 vssd1 vccd1 vccd1 _16617_/A0 sky130_fd_sc_hd__buf_2
X_09879_ _18534_/Q _18409_/Q _10054_/S vssd1 vssd1 vccd1 vccd1 _09879_/X sky130_fd_sc_hd__mux2_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _18564_/Q _11663_/A _11706_/B _11732_/Y vssd1 vssd1 vccd1 vccd1 _11910_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _13135_/S _12875_/X _12880_/X _13194_/S vssd1 vssd1 vccd1 vccd1 _12890_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_302 _18112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 _18116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 _18109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11841_ _11841_/A _11864_/B vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__or2_2
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_335 _14663_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 _10364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_357 _12461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_368 _16110_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11772_ _11799_/A _15039_/B _11726_/B vssd1 vssd1 vccd1 vccd1 _11772_/X sky130_fd_sc_hd__a21o_1
XFILLER_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14560_ _14586_/A _14560_/B vssd1 vssd1 vccd1 vccd1 _18388_/D sky130_fd_sc_hd__or2_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_379 _14940_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10723_ _18070_/Q _10816_/A2 _10722_/X _10719_/S vssd1 vssd1 vccd1 vccd1 _10723_/X
+ sky130_fd_sc_hd__o211a_1
X_13511_ _13545_/A _13511_/B vssd1 vssd1 vccd1 vccd1 _13511_/Y sky130_fd_sc_hd__nand2_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14491_ _16593_/A0 _18341_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _18341_/D sky130_fd_sc_hd__mux2_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _16594_/A0 _18845_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _18845_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10654_ _10881_/S1 _10643_/X _10653_/X _11621_/C1 vssd1 vssd1 vccd1 vccd1 _10654_/X
+ sky130_fd_sc_hd__o211a_1
X_13442_ _13937_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13442_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13373_ _19406_/Q _12579_/Y _12771_/X _13372_/X _12581_/Y vssd1 vssd1 vccd1 vccd1
+ _13373_/X sky130_fd_sc_hd__a221o_1
X_16161_ _17625_/A _16260_/B vssd1 vssd1 vccd1 vccd1 _16161_/Y sky130_fd_sc_hd__nand2_2
XFILLER_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10585_ _10581_/X _10582_/X _10668_/S vssd1 vssd1 vccd1 vccd1 _10585_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15112_ _15112_/A _15112_/B vssd1 vssd1 vccd1 vccd1 _15112_/Y sky130_fd_sc_hd__nor2_4
XFILLER_182_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12324_ _08932_/A _08912_/Y _08927_/Y _17793_/Q _08942_/B vssd1 vssd1 vccd1 vccd1
+ _12324_/Y sky130_fd_sc_hd__o2111ai_1
X_16092_ _16096_/A1 _16091_/Y _17725_/C1 vssd1 vssd1 vccd1 vccd1 _18748_/D sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_1_wb_clk_i _19652_/A vssd1 vssd1 vccd1 vccd1 _19637_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_181_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12255_ _17884_/Q _12251_/B _12254_/Y vssd1 vssd1 vccd1 vccd1 _17884_/D sky130_fd_sc_hd__o21a_1
X_15043_ _17342_/A _15043_/B _15043_/C vssd1 vssd1 vccd1 vccd1 _18530_/D sky130_fd_sc_hd__and3_1
XFILLER_253_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11206_ _11616_/S _11205_/X _11508_/B1 vssd1 vssd1 vccd1 vccd1 _11206_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12186_ _17859_/Q _12186_/B vssd1 vssd1 vccd1 vccd1 _12192_/C sky130_fd_sc_hd__and2_2
XFILLER_269_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18802_ _19644_/CLK _18802_/D vssd1 vssd1 vccd1 vccd1 _18802_/Q sky130_fd_sc_hd__dfxtp_1
X_11137_ _11138_/A _11138_/B vssd1 vssd1 vccd1 vccd1 _13487_/S sky130_fd_sc_hd__and2_4
XFILLER_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16994_ _17569_/A _17044_/A2 _16993_/X _17322_/A vssd1 vssd1 vccd1 vccd1 _19333_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18733_ _18734_/CLK _18733_/D vssd1 vssd1 vccd1 vccd1 _18733_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_283_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15945_ _18690_/Q _15948_/A2 _15923_/C _15944_/X _15945_/C1 vssd1 vssd1 vccd1 vccd1
+ _15945_/X sky130_fd_sc_hd__a221o_1
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11068_ _18988_/Q _11300_/B vssd1 vssd1 vccd1 vccd1 _11068_/X sky130_fd_sc_hd__or2_1
XFILLER_83_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10019_ _11566_/A1 _18133_/Q _18779_/Q _11581_/S _12320_/A vssd1 vssd1 vccd1 vccd1
+ _10020_/C sky130_fd_sc_hd__a221o_1
X_18664_ _18666_/CLK _18664_/D vssd1 vssd1 vccd1 vccd1 _18664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15876_ _18667_/Q _15853_/Y _15906_/B1 vssd1 vssd1 vccd1 vccd1 _15876_/X sky130_fd_sc_hd__a21o_1
XFILLER_236_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _19488_/Q _15088_/X _17556_/A _17202_/B _17556_/X vssd1 vssd1 vccd1 vccd1
+ _17615_/X sky130_fd_sc_hd__a221o_1
XFILLER_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14827_ _14823_/Y _14826_/X _14950_/B1 vssd1 vssd1 vccd1 vccd1 _14827_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18595_ _19619_/CLK _18595_/D vssd1 vssd1 vccd1 vccd1 _18595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_252_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17546_ _18131_/Q _17546_/A2 _17219_/A _17545_/X vssd1 vssd1 vccd1 vccd1 _17546_/X
+ sky130_fd_sc_hd__o211a_1
X_14758_ _18477_/Q _14720_/A _14757_/Y _12243_/A vssd1 vssd1 vccd1 vccd1 _18477_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_251_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13709_ _09777_/A _12762_/A _13808_/C1 _13708_/Y vssd1 vssd1 vccd1 vccd1 _13709_/X
+ sky130_fd_sc_hd__a211o_4
X_17477_ _18118_/Q _17539_/C1 _17475_/X _17476_/X vssd1 vssd1 vccd1 vccd1 _17477_/X
+ sky130_fd_sc_hd__a22o_1
X_14689_ _14417_/C _14692_/A2 _12276_/B vssd1 vssd1 vccd1 vccd1 _14689_/Y sky130_fd_sc_hd__a21oi_1
X_19216_ _19216_/CLK _19216_/D vssd1 vssd1 vccd1 vccd1 _19216_/Q sky130_fd_sc_hd__dfxtp_1
X_16428_ _19036_/Q _16593_/A0 _16457_/S vssd1 vssd1 vccd1 vccd1 _19036_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19147_ _19147_/CLK _19147_/D vssd1 vssd1 vccd1 vccd1 _19147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16359_ _16359_/A _16459_/C vssd1 vssd1 vccd1 vccd1 _16359_/X sky130_fd_sc_hd__or2_4
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19078_ _19140_/CLK _19078_/D vssd1 vssd1 vccd1 vccd1 _19078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18029_ _19599_/CLK _18029_/D vssd1 vssd1 vccd1 vccd1 _18029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_278_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09802_ _18629_/Q _11617_/S vssd1 vssd1 vccd1 vccd1 _09802_/X sky130_fd_sc_hd__or2_1
XFILLER_87_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09733_ _09735_/A _12609_/B vssd1 vssd1 vccd1 vccd1 _12999_/S sky130_fd_sc_hd__nand2_4
XFILLER_68_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09664_ _10262_/A1 _18137_/Q _18783_/Q _09671_/S _11397_/A1 vssd1 vssd1 vccd1 vccd1
+ _09664_/X sky130_fd_sc_hd__a221o_1
XFILLER_28_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09595_ _09593_/X _09594_/X _09718_/S vssd1 vssd1 vccd1 vccd1 _09595_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_71_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19565_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ _19645_/Q _18934_/Q _10370_/S vssd1 vssd1 vccd1 vccd1 _10370_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09029_ _17921_/Q _09031_/S vssd1 vssd1 vccd1 vccd1 _09902_/B sky130_fd_sc_hd__nand2_2
XFILLER_152_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _17895_/Q _12052_/A2 _12039_/X _13100_/A vssd1 vssd1 vccd1 vccd1 _17797_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1704 _09086_/A vssd1 vssd1 vccd1 vccd1 _11588_/B1 sky130_fd_sc_hd__clkbuf_16
Xfanout1715 _12492_/A vssd1 vssd1 vccd1 vccd1 _16848_/S sky130_fd_sc_hd__buf_8
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1726 _08828_/A vssd1 vssd1 vccd1 vccd1 _16821_/A sky130_fd_sc_hd__buf_6
Xfanout1737 _18339_/Q vssd1 vssd1 vccd1 vccd1 _09655_/S sky130_fd_sc_hd__buf_6
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout750 _13046_/A1 vssd1 vssd1 vccd1 vccd1 _13414_/A sky130_fd_sc_hd__clkbuf_4
Xfanout1748 _18105_/Q vssd1 vssd1 vccd1 vccd1 _14214_/A sky130_fd_sc_hd__buf_12
XFILLER_77_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout761 _17670_/A0 vssd1 vssd1 vccd1 vccd1 _17703_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout1759 _09099_/A vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__buf_12
XFILLER_265_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout772 _17658_/Y vssd1 vssd1 vccd1 vccd1 _17687_/S sky130_fd_sc_hd__buf_12
X_13991_ _17960_/Q _14034_/B _13990_/Y _14001_/C1 vssd1 vssd1 vccd1 vccd1 _17960_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout783 _16590_/S vssd1 vssd1 vccd1 vccd1 _16586_/S sky130_fd_sc_hd__buf_12
XFILLER_218_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout794 _16326_/Y vssd1 vssd1 vccd1 vccd1 _16352_/S sky130_fd_sc_hd__clkbuf_16
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _18590_/Q _15746_/C vssd1 vssd1 vccd1 vccd1 _15730_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _12793_/X _12805_/X _12942_/S vssd1 vssd1 vccd1 vccd1 _12942_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _19449_/Q _15661_/B vssd1 vssd1 vccd1 vccd1 _15661_/X sky130_fd_sc_hd__or2_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12873_ _12942_/S _12670_/X _12872_/Y vssd1 vssd1 vccd1 vccd1 _12873_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_110 _11751_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_121 _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_132 _11814_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _19491_/Q _17462_/B _17399_/X vssd1 vssd1 vccd1 vccd1 _19491_/D sky130_fd_sc_hd__o21ba_1
X_14612_ _17671_/A0 _18419_/Q _14628_/S vssd1 vssd1 vccd1 vccd1 _18419_/D sky130_fd_sc_hd__mux2_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _11857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18380_ _19483_/CLK _18380_/D vssd1 vssd1 vccd1 vccd1 _18380_/Q sky130_fd_sc_hd__dfxtp_4
X_11824_ _11824_/A _11858_/B vssd1 vssd1 vccd1 vccd1 _11827_/B sky130_fd_sc_hd__or2_2
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _19477_/Q _15591_/Y _15781_/S vssd1 vssd1 vccd1 vccd1 _15592_/X sky130_fd_sc_hd__mux2_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _11872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_165 _12949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_176 _14002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_187 _13677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17331_ _19463_/Q _17573_/A _17377_/S vssd1 vssd1 vccd1 vccd1 _17332_/B sky130_fd_sc_hd__mux2_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _18380_/Q _14559_/A2 _14559_/B1 input39/X vssd1 vssd1 vccd1 vccd1 _14544_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_198 _13886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _18573_/Q _14522_/A2 _11818_/B _13258_/A vssd1 vssd1 vccd1 vccd1 _11755_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17262_ _19438_/Q _17310_/B vssd1 vssd1 vccd1 vccd1 _17262_/Y sky130_fd_sc_hd__nand2_1
X_10706_ _10704_/X _10705_/X _10706_/S vssd1 vssd1 vccd1 vccd1 _10707_/B sky130_fd_sc_hd__mux2_1
X_14474_ _18326_/Q _16611_/A0 _14486_/S vssd1 vssd1 vccd1 vccd1 _18326_/D sky130_fd_sc_hd__mux2_1
X_11686_ _11686_/A _13622_/B _13611_/B _11686_/D vssd1 vssd1 vccd1 vccd1 _11686_/X
+ sky130_fd_sc_hd__or4_1
X_19001_ _19225_/CLK _19001_/D vssd1 vssd1 vccd1 vccd1 _19001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16213_ _17710_/A0 _18829_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _18829_/D sky130_fd_sc_hd__mux2_1
X_13425_ _19247_/Q _13425_/A2 _13425_/B1 _19279_/Q vssd1 vssd1 vccd1 vccd1 _13425_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10637_ _10623_/A _10636_/Y _10623_/Y _11333_/A1 vssd1 vssd1 vccd1 vccd1 _10637_/Y
+ sky130_fd_sc_hd__o211ai_2
X_17193_ _17214_/A _17193_/B vssd1 vssd1 vccd1 vccd1 _17513_/A sky130_fd_sc_hd__nand2_2
XFILLER_127_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16144_ _18725_/Q _18724_/Q vssd1 vssd1 vccd1 vccd1 _16145_/C sky130_fd_sc_hd__nor2_1
XFILLER_155_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13356_ _12739_/S _12896_/Y _13355_/X vssd1 vssd1 vccd1 vccd1 _13356_/X sky130_fd_sc_hd__a21o_1
X_10568_ _10566_/X _10567_/X _10643_/S vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12307_ _16819_/B vssd1 vssd1 vccd1 vccd1 _14934_/D sky130_fd_sc_hd__inv_2
XFILLER_6_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16075_ _16075_/A _16075_/B _16075_/C vssd1 vssd1 vccd1 vccd1 _16075_/Y sky130_fd_sc_hd__nand3_1
X_10499_ _10033_/S _10498_/X _10497_/X _11274_/S1 vssd1 vssd1 vccd1 vccd1 _10499_/X
+ sky130_fd_sc_hd__a211o_1
X_13287_ _13757_/A _13996_/B _13274_/Y vssd1 vssd1 vccd1 vccd1 _13287_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15026_ _18515_/Q input192/X _15038_/S vssd1 vssd1 vccd1 vccd1 _18515_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12238_ _17878_/Q _12240_/C _12237_/Y vssd1 vssd1 vccd1 vccd1 _17878_/D sky130_fd_sc_hd__o21a_1
XFILLER_130_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12169_ _16811_/A _12169_/B _12170_/B vssd1 vssd1 vccd1 vccd1 _17852_/D sky130_fd_sc_hd__nor3_1
XFILLER_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16977_ _17051_/A _16977_/B vssd1 vssd1 vccd1 vccd1 _17591_/C sky130_fd_sc_hd__nand2_8
XFILLER_232_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput5 coreIndex[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_6
XFILLER_65_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15928_ _18685_/Q _15943_/A2 _15927_/X _15946_/C1 vssd1 vssd1 vccd1 vccd1 _18685_/D
+ sky130_fd_sc_hd__o211a_1
X_18716_ _19142_/CLK _18716_/D vssd1 vssd1 vccd1 vccd1 _18716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_283_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18647_ _19586_/CLK _18647_/D vssd1 vssd1 vccd1 vccd1 _18647_/Q sky130_fd_sc_hd__dfxtp_4
X_15859_ _18662_/Q _15949_/A2 _15857_/X _15858_/X _14205_/A vssd1 vssd1 vccd1 vccd1
+ _18662_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09380_ _19626_/Q _18915_/Q _10141_/S vssd1 vssd1 vccd1 vccd1 _09380_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18578_ _19506_/CLK _18578_/D vssd1 vssd1 vccd1 vccd1 _18578_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_252_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17529_ _17202_/Y _17517_/B _17527_/X _17528_/Y _17285_/A vssd1 vssd1 vccd1 vccd1
+ _17529_/X sky130_fd_sc_hd__a41o_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput320 _11767_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[23] sky130_fd_sc_hd__buf_4
XFILLER_273_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput331 _11749_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[8] sky130_fd_sc_hd__buf_4
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput342 _11844_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[17] sky130_fd_sc_hd__buf_4
XFILLER_126_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput353 _11890_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[27] sky130_fd_sc_hd__buf_4
XFILLER_0_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput364 _11806_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[8] sky130_fd_sc_hd__buf_4
XFILLER_102_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput375 _14487_/B vssd1 vssd1 vccd1 vccd1 csb1[1] sky130_fd_sc_hd__buf_4
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput386 _11939_/X vssd1 vssd1 vccd1 vccd1 din0[19] sky130_fd_sc_hd__buf_4
Xoutput397 _11949_/X vssd1 vssd1 vccd1 vccd1 din0[29] sky130_fd_sc_hd__buf_4
XFILLER_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09716_ _18311_/Q _17762_/Q _09724_/S vssd1 vssd1 vccd1 vccd1 _09716_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09647_ _12614_/B _09647_/B vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__xor2_4
XFILLER_216_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09578_ _19040_/Q _19008_/Q _10362_/S vssd1 vssd1 vccd1 vccd1 _09578_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ _11541_/A _10754_/A _11541_/B vssd1 vssd1 vccd1 vccd1 _11540_/X sky130_fd_sc_hd__o21ba_1
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11471_ _19047_/Q _19015_/Q _11481_/C vssd1 vssd1 vccd1 vccd1 _11471_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ _18652_/Q _10424_/S vssd1 vssd1 vccd1 vccd1 _10422_/X sky130_fd_sc_hd__or2_1
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13210_ _19401_/Q _12570_/A _13244_/B1 vssd1 vssd1 vccd1 vccd1 _13210_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ _18706_/Q _18093_/Q _14200_/S vssd1 vssd1 vccd1 vccd1 _14191_/B sky130_fd_sc_hd__mux2_1
XFILLER_136_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10353_ _19094_/Q _18998_/Q _10353_/S vssd1 vssd1 vccd1 vccd1 _10353_/X sky130_fd_sc_hd__mux2_1
X_13141_ _11745_/A _13316_/B _12836_/Y _13127_/A _13260_/A vssd1 vssd1 vccd1 vccd1
+ _13141_/Y sky130_fd_sc_hd__a221oi_4
XFILLER_152_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13072_ _15875_/A _12506_/X _13060_/X _13071_/X _12510_/X vssd1 vssd1 vccd1 vccd1
+ _13072_/X sky130_fd_sc_hd__o221a_1
XFILLER_152_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10284_ _10275_/S _10277_/X _10276_/X _09429_/S vssd1 vssd1 vccd1 vccd1 _10284_/X
+ sky130_fd_sc_hd__a211o_1
X_16900_ _16960_/A _16900_/B vssd1 vssd1 vccd1 vccd1 _19309_/D sky130_fd_sc_hd__and2_1
X_12023_ _12023_/A _12433_/B vssd1 vssd1 vccd1 vccd1 _12023_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1501 _09498_/S vssd1 vssd1 vccd1 vccd1 _09724_/S sky130_fd_sc_hd__buf_4
XFILLER_105_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17880_ _19324_/CLK _17880_/D vssd1 vssd1 vccd1 vccd1 _17880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1512 _10199_/S vssd1 vssd1 vccd1 vccd1 _10348_/S sky130_fd_sc_hd__clkbuf_8
Xfanout1523 fanout1524/X vssd1 vssd1 vccd1 vccd1 _10426_/S sky130_fd_sc_hd__buf_4
XFILLER_250_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1534 _10653_/A1 vssd1 vssd1 vccd1 vccd1 _10275_/S sky130_fd_sc_hd__buf_8
XFILLER_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16831_ _16831_/A _16831_/B vssd1 vssd1 vccd1 vccd1 _17052_/A sky130_fd_sc_hd__nand2_1
Xfanout1545 _08899_/Y vssd1 vssd1 vccd1 vccd1 _10649_/A1 sky130_fd_sc_hd__buf_4
Xfanout1556 _09381_/S vssd1 vssd1 vccd1 vccd1 _10205_/S sky130_fd_sc_hd__buf_6
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1567 _11508_/B1 vssd1 vssd1 vccd1 vccd1 _11279_/B1 sky130_fd_sc_hd__clkbuf_16
Xfanout1578 _11507_/S vssd1 vssd1 vccd1 vccd1 _11514_/S sky130_fd_sc_hd__buf_8
XFILLER_219_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout580 _12338_/Y vssd1 vssd1 vccd1 vccd1 _12421_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_120_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1589 _10211_/A1 vssd1 vssd1 vccd1 vccd1 _11046_/S1 sky130_fd_sc_hd__buf_8
Xfanout591 _12023_/Y vssd1 vssd1 vccd1 vccd1 _12073_/B sky130_fd_sc_hd__buf_4
X_19550_ _19553_/CLK _19550_/D vssd1 vssd1 vccd1 vccd1 _19550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16762_ _19274_/Q _16762_/B vssd1 vssd1 vccd1 vccd1 _16767_/C sky130_fd_sc_hd__and2_2
XFILLER_265_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13974_ _17952_/Q _14028_/A vssd1 vssd1 vccd1 vccd1 _13974_/X sky130_fd_sc_hd__or2_1
XFILLER_76_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18501_ _18501_/CLK _18501_/D vssd1 vssd1 vccd1 vccd1 _18501_/Q sky130_fd_sc_hd__dfxtp_1
X_15713_ _15713_/A _15713_/B vssd1 vssd1 vccd1 vccd1 _15715_/A sky130_fd_sc_hd__nand2_1
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19481_ _19481_/CLK _19481_/D vssd1 vssd1 vccd1 vccd1 _19481_/Q sky130_fd_sc_hd__dfxtp_2
X_12925_ _18102_/Q _12788_/B _18104_/Q _18103_/Q vssd1 vssd1 vccd1 vccd1 _13028_/C
+ sky130_fd_sc_hd__o211a_4
X_16693_ _19250_/Q _16699_/D _16692_/Y vssd1 vssd1 vccd1 vccd1 _19250_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18432_ _19092_/CLK _18432_/D vssd1 vssd1 vccd1 vccd1 _18432_/Q sky130_fd_sc_hd__dfxtp_1
X_15644_ _15686_/A _15644_/B vssd1 vssd1 vccd1 vccd1 _15645_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _19362_/Q _12516_/Y _12849_/X _12855_/X vssd1 vssd1 vccd1 vccd1 _12856_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_261_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18363_ _19641_/CLK _18363_/D vssd1 vssd1 vccd1 vccd1 _18363_/Q sky130_fd_sc_hd__dfxtp_1
X_11807_ _11820_/A _11807_/B vssd1 vssd1 vccd1 vccd1 _11807_/Y sky130_fd_sc_hd__nor2_2
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15575_ _18122_/Q _15763_/A2 _15574_/X _15481_/B vssd1 vssd1 vccd1 vccd1 _15639_/A
+ sky130_fd_sc_hd__o22a_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12787_ _18102_/Q _12788_/B vssd1 vssd1 vccd1 vccd1 _12868_/B sky130_fd_sc_hd__nor2_2
XFILLER_221_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _14268_/A _17214_/A _17214_/Y _17313_/B vssd1 vssd1 vccd1 vccd1 _17314_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_203_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ input9/X _14528_/B vssd1 vssd1 vccd1 vccd1 _14527_/B sky130_fd_sc_hd__nor2_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18294_ _18593_/CLK _18294_/D vssd1 vssd1 vccd1 vccd1 _18294_/Q sky130_fd_sc_hd__dfxtp_1
X_11738_ _18566_/Q _11741_/A2 _11769_/B1 _11737_/X vssd1 vssd1 vccd1 vccd1 _11738_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17245_ _18109_/Q _17129_/A _17433_/A _17244_/B vssd1 vssd1 vccd1 vccd1 _17245_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_186_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14457_ _18309_/Q _17694_/A0 _14477_/S vssd1 vssd1 vccd1 vccd1 _18309_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11669_ _12638_/A _11669_/B vssd1 vssd1 vccd1 vccd1 _13676_/B sky130_fd_sc_hd__xnor2_4
XFILLER_174_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13408_ _13408_/A vssd1 vssd1 vccd1 vccd1 _13408_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17176_ _19410_/Q fanout536/X _17483_/A _17120_/B vssd1 vssd1 vccd1 vccd1 _17177_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_128_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14388_ _17695_/A0 _18239_/Q _14416_/S vssd1 vssd1 vccd1 vccd1 _18239_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16127_ _18766_/Q _16139_/B vssd1 vssd1 vccd1 vccd1 _16127_/Y sky130_fd_sc_hd__nand2_1
X_13339_ _19469_/Q _12529_/Y _12578_/Y _19341_/Q _13338_/X vssd1 vssd1 vccd1 vccd1
+ _13339_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16058_ _16063_/B _16055_/A _16057_/X _16039_/X vssd1 vssd1 vccd1 vccd1 _16058_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15009_ _15009_/A1 _18272_/Q _15008_/Y input205/X vssd1 vssd1 vccd1 vccd1 _15009_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_69_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08880_ _12323_/A _09073_/D _12320_/C _08880_/D vssd1 vssd1 vccd1 vccd1 _08882_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_285_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09501_ _12962_/A0 _09499_/X _09500_/X _08895_/A vssd1 vssd1 vccd1 vccd1 _09501_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_271_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09432_ _08904_/A _09411_/Y _09417_/Y _09424_/Y _09431_/X vssd1 vssd1 vccd1 vccd1
+ _09432_/X sky130_fd_sc_hd__o32a_4
XFILLER_213_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09363_ _11024_/A1 _09362_/X _11023_/B1 vssd1 vssd1 vccd1 vccd1 _09363_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09294_ _19627_/Q _18916_/Q _09302_/S vssd1 vssd1 vccd1 vccd1 _09294_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_10 _18528_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _14980_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_32 _17073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 _12600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_54 _09743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_87 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_98 _11067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10971_ _11360_/A1 _19605_/Q _19573_/Q _11340_/B2 vssd1 vssd1 vccd1 vccd1 _10971_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12710_ _12705_/X _12709_/X _12878_/S vssd1 vssd1 vccd1 vccd1 _12710_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13690_ _17846_/Q _13846_/B _13683_/X _13689_/X vssd1 vssd1 vccd1 vccd1 _13690_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12641_ _12641_/A _12641_/B vssd1 vssd1 vccd1 vccd1 _13615_/B sky130_fd_sc_hd__or2_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15360_ _12665_/A _12318_/A _15437_/B1 _15330_/B _15361_/B vssd1 vssd1 vccd1 vccd1
+ _15385_/A sky130_fd_sc_hd__a2111o_1
X_12572_ _12572_/A _12572_/B _12572_/C _12503_/Y vssd1 vssd1 vccd1 vccd1 _12584_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14311_ _18168_/Q _16595_/A0 _14325_/S vssd1 vssd1 vccd1 vccd1 _18168_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11523_ _13316_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _13311_/A sky130_fd_sc_hd__nor2_4
X_15291_ _15262_/A _15262_/B _15268_/Y vssd1 vssd1 vccd1 vccd1 _15293_/B sky130_fd_sc_hd__o21a_1
XFILLER_200_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17030_ _17190_/B _17046_/A2 _17029_/X _17106_/C1 vssd1 vssd1 vccd1 vccd1 _19351_/D
+ sky130_fd_sc_hd__o211a_1
X_14242_ _18119_/Q _14244_/B vssd1 vssd1 vccd1 vccd1 _14242_/X sky130_fd_sc_hd__or2_1
X_11454_ _19079_/Q _11455_/S _11453_/X _11464_/C1 vssd1 vssd1 vccd1 vccd1 _11454_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ _09135_/S _10400_/X _10404_/X vssd1 vssd1 vccd1 vccd1 _10405_/X sky130_fd_sc_hd__o21a_1
XFILLER_139_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11385_ _18420_/Q _10101_/B _11384_/X _10403_/S vssd1 vssd1 vccd1 vccd1 _11385_/X
+ sky130_fd_sc_hd__o211a_1
X_14173_ _16968_/A _14173_/B vssd1 vssd1 vccd1 vccd1 _18084_/D sky130_fd_sc_hd__and2_1
XFILLER_183_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13124_ _13936_/B2 _13122_/Y _13123_/X _13185_/A vssd1 vssd1 vccd1 vccd1 _13124_/X
+ sky130_fd_sc_hd__a211o_1
X_10336_ _10336_/A _10336_/B vssd1 vssd1 vccd1 vccd1 _10336_/X sky130_fd_sc_hd__or2_2
XFILLER_194_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18981_ _19564_/CLK _18981_/D vssd1 vssd1 vccd1 vccd1 _18981_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17932_ _18627_/CLK _17932_/D vssd1 vssd1 vccd1 vccd1 _17932_/Q sky130_fd_sc_hd__dfxtp_2
X_10267_ _09463_/S _10266_/X _10996_/B1 vssd1 vssd1 vccd1 vccd1 _10267_/X sky130_fd_sc_hd__o21a_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _18107_/Q _13055_/B vssd1 vssd1 vccd1 vccd1 _13056_/B sky130_fd_sc_hd__nor2_1
XFILLER_279_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1320 _09106_/B vssd1 vssd1 vccd1 vccd1 _11570_/B1 sky130_fd_sc_hd__buf_8
XFILLER_266_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12006_ _17773_/Q _17674_/A0 _12013_/S vssd1 vssd1 vccd1 vccd1 _17773_/D sky130_fd_sc_hd__mux2_1
X_17863_ _17865_/CLK _17863_/D vssd1 vssd1 vccd1 vccd1 _17863_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1331 _10004_/A1 vssd1 vssd1 vccd1 vccd1 _10707_/A sky130_fd_sc_hd__buf_6
X_10198_ _18336_/Q _17787_/Q _10206_/S vssd1 vssd1 vccd1 vccd1 _10198_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1342 _10618_/S vssd1 vssd1 vccd1 vccd1 _10930_/S sky130_fd_sc_hd__buf_4
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1353 _09914_/C1 vssd1 vssd1 vccd1 vccd1 _09135_/S sky130_fd_sc_hd__buf_6
XFILLER_93_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1364 _11325_/S vssd1 vssd1 vccd1 vccd1 _10864_/S sky130_fd_sc_hd__buf_6
X_19602_ _19602_/CLK _19602_/D vssd1 vssd1 vccd1 vccd1 _19602_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1375 _10634_/S0 vssd1 vssd1 vccd1 vccd1 _09108_/B sky130_fd_sc_hd__buf_6
XFILLER_282_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16814_ _19293_/Q _19292_/Q _16810_/B _19294_/Q vssd1 vssd1 vccd1 vccd1 _16816_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_281_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17794_ _19650_/CLK _17794_/D vssd1 vssd1 vccd1 vccd1 _17794_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1386 _09843_/S vssd1 vssd1 vccd1 vccd1 fanout1386/X sky130_fd_sc_hd__buf_4
Xfanout1397 _10249_/S vssd1 vssd1 vccd1 vccd1 _10253_/C sky130_fd_sc_hd__buf_6
X_16745_ _19268_/Q _16746_/B vssd1 vssd1 vccd1 vccd1 _16747_/B sky130_fd_sc_hd__nor2_1
XFILLER_235_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19533_ _19533_/CLK _19533_/D vssd1 vssd1 vccd1 vccd1 _19533_/Q sky130_fd_sc_hd__dfxtp_1
X_13957_ _13931_/A _13955_/X _13956_/Y _13958_/A _13294_/A vssd1 vssd1 vccd1 vccd1
+ _13957_/X sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_199_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19607_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_250_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12908_ _19235_/Q _13495_/A2 _13495_/B1 _19267_/Q vssd1 vssd1 vccd1 vccd1 _12908_/X
+ sky130_fd_sc_hd__a22o_1
X_19464_ _19464_/CLK _19464_/D vssd1 vssd1 vccd1 vccd1 _19464_/Q sky130_fd_sc_hd__dfxtp_2
X_16676_ _19247_/Q _19246_/Q _19245_/Q vssd1 vssd1 vccd1 vccd1 _16677_/D sky130_fd_sc_hd__and3_1
XFILLER_234_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13888_ _13930_/A1 _13874_/X _13930_/B1 vssd1 vssd1 vccd1 vccd1 _13888_/X sky130_fd_sc_hd__o21a_1
XFILLER_146_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_128_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19229_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18415_ _19075_/CLK _18415_/D vssd1 vssd1 vccd1 vccd1 _18415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15627_ _15610_/B _15612_/B _15610_/A vssd1 vssd1 vccd1 vccd1 _15631_/A sky130_fd_sc_hd__o21bai_2
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12839_ _12878_/S _09984_/B _13912_/B1 _12838_/X vssd1 vssd1 vccd1 vccd1 _12839_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19395_ _19525_/CLK _19395_/D vssd1 vssd1 vccd1 vccd1 _19395_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18346_ _18445_/CLK _18346_/D vssd1 vssd1 vccd1 vccd1 _18346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15558_ _15558_/A _15558_/B vssd1 vssd1 vccd1 vccd1 _15558_/X sky130_fd_sc_hd__or2_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14509_ _17678_/A0 _18359_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _18359_/D sky130_fd_sc_hd__mux2_1
X_18277_ _18279_/CLK _18277_/D vssd1 vssd1 vccd1 vccd1 _18277_/Q sky130_fd_sc_hd__dfxtp_1
X_15489_ _15557_/B _15489_/B vssd1 vssd1 vccd1 vccd1 _15489_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_163_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17228_ _17226_/Y _17227_/X _17141_/A vssd1 vssd1 vccd1 vccd1 _19426_/D sky130_fd_sc_hd__a21oi_1
XFILLER_190_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput30 core_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput41 core_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
Xinput52 dout0[18] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput63 dout0[28] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17159_ _17159_/A _17159_/B vssd1 vssd1 vccd1 vccd1 _19404_/D sky130_fd_sc_hd__nor2_1
XFILLER_7_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput74 dout0[38] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_2
Xinput85 dout0[48] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_2
Xinput96 dout0[58] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09981_ _09948_/B _09980_/Y _09948_/X vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__a21boi_4
XFILLER_171_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08932_ _08932_/A _12051_/A _17802_/Q _12053_/A vssd1 vssd1 vccd1 vccd1 _08932_/X
+ sky130_fd_sc_hd__or4bb_1
XFILLER_103_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08863_ _11689_/A vssd1 vssd1 vccd1 vccd1 _08863_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09415_ _18850_/Q _18882_/Q _19042_/Q _19010_/Q _09428_/B2 _11199_/S1 vssd1 vssd1
+ vccd1 vccd1 _09415_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09346_ _10169_/S _09344_/X _09345_/X vssd1 vssd1 vccd1 vccd1 _09346_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09277_ _11024_/A1 _09276_/X _11257_/C1 vssd1 vssd1 vccd1 vccd1 _09277_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11170_ _09845_/S _11169_/X _10689_/S vssd1 vssd1 vccd1 vccd1 _11170_/X sky130_fd_sc_hd__a21o_1
XFILLER_162_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10121_ _11488_/A _10121_/B vssd1 vssd1 vccd1 vccd1 _10121_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10052_ _19099_/Q _19131_/Q _10054_/S vssd1 vssd1 vccd1 vccd1 _10052_/X sky130_fd_sc_hd__mux2_1
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860_ _18487_/Q _15001_/A2 _14859_/Y _16808_/A vssd1 vssd1 vccd1 vccd1 _18487_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _11639_/A _13794_/B _12648_/X vssd1 vssd1 vccd1 vccd1 _13812_/B sky130_fd_sc_hd__a21o_2
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14791_ _14789_/X _14790_/X _14964_/B1 vssd1 vssd1 vccd1 vccd1 _14791_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16530_ _16530_/A0 _19135_/Q _16554_/S vssd1 vssd1 vccd1 vccd1 _19135_/D sky130_fd_sc_hd__mux2_1
X_13742_ _17944_/Q _13742_/A2 _13741_/X _14179_/A vssd1 vssd1 vccd1 vccd1 _17944_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_232_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10954_ _11352_/A1 _18613_/Q _18184_/Q _11353_/B2 vssd1 vssd1 vccd1 vccd1 _10954_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16461_ _16461_/A0 _19068_/Q _16488_/S vssd1 vssd1 vccd1 vccd1 _19068_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13673_ _18123_/Q _13704_/C vssd1 vssd1 vccd1 vccd1 _13673_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10885_ _10883_/X _10884_/X _11127_/S vssd1 vssd1 vccd1 vccd1 _10885_/X sky130_fd_sc_hd__mux2_1
XFILLER_231_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18200_ _18817_/CLK _18200_/D vssd1 vssd1 vccd1 vccd1 _18200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15412_ _18576_/Q _15412_/B vssd1 vssd1 vccd1 vccd1 _15465_/C sky130_fd_sc_hd__and2_2
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19180_ _19621_/CLK _19180_/D vssd1 vssd1 vccd1 vccd1 _19180_/Q sky130_fd_sc_hd__dfxtp_1
X_12624_ _12624_/A _12624_/B vssd1 vssd1 vccd1 vccd1 _13311_/B sky130_fd_sc_hd__nand2_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16392_ _17800_/Q _16392_/B _16392_/C vssd1 vssd1 vccd1 vccd1 _16591_/B sky130_fd_sc_hd__and3_2
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18131_ _18593_/CLK _18131_/D vssd1 vssd1 vccd1 vccd1 _18131_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15343_ _15388_/C _15342_/Y _15124_/X vssd1 vssd1 vccd1 vccd1 _15343_/Y sky130_fd_sc_hd__o21ai_1
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ _12575_/A _12561_/B vssd1 vssd1 vccd1 vccd1 _12555_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ _11506_/A1 _19111_/Q _19143_/Q _10424_/S vssd1 vssd1 vccd1 vccd1 _11506_/X
+ sky130_fd_sc_hd__a22o_1
X_18062_ _19226_/CLK _18062_/D vssd1 vssd1 vccd1 vccd1 _18062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15274_ _17166_/A _15274_/B _15274_/C vssd1 vssd1 vccd1 vccd1 _15274_/X sky130_fd_sc_hd__and3_1
XFILLER_129_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12486_ _12492_/A _12486_/B vssd1 vssd1 vccd1 vccd1 _12486_/X sky130_fd_sc_hd__and2_1
XFILLER_184_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17013_ _19343_/Q _17045_/B vssd1 vssd1 vccd1 vccd1 _17013_/X sky130_fd_sc_hd__or2_1
X_14225_ _18284_/Q _14224_/B _14224_/Y _17352_/A vssd1 vssd1 vccd1 vccd1 _18110_/D
+ sky130_fd_sc_hd__o211a_1
X_11437_ _11428_/A _11436_/X _11515_/B1 vssd1 vssd1 vccd1 vccd1 _11437_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14156_ _14156_/A0 _13316_/B _14156_/S vssd1 vssd1 vccd1 vccd1 _14156_/X sky130_fd_sc_hd__mux2_1
X_11368_ _11368_/A _12596_/B vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__and2_2
XFILLER_180_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13107_ _19529_/Q _13372_/S vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__or2_1
X_10319_ _18263_/Q _18838_/Q _10687_/S vssd1 vssd1 vccd1 vccd1 _10319_/X sky130_fd_sc_hd__mux2_1
X_14087_ _17703_/A0 _18027_/Q _14106_/S vssd1 vssd1 vccd1 vccd1 _18027_/D sky130_fd_sc_hd__mux2_1
X_18964_ _19620_/CLK _18964_/D vssd1 vssd1 vccd1 vccd1 _18964_/Q sky130_fd_sc_hd__dfxtp_1
X_11299_ _17934_/Q _08946_/Y _11298_/X _11451_/B2 vssd1 vssd1 vccd1 vccd1 _11299_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17915_ _18881_/CLK _17915_/D vssd1 vssd1 vccd1 vccd1 _17915_/Q sky130_fd_sc_hd__dfxtp_4
X_13038_ _13354_/A _13038_/B vssd1 vssd1 vccd1 vccd1 _13038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18895_ _19055_/CLK _18895_/D vssd1 vssd1 vccd1 vccd1 _18895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1150 _13916_/A vssd1 vssd1 vccd1 vccd1 _13294_/A sky130_fd_sc_hd__buf_6
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1161 _16003_/A2 vssd1 vssd1 vccd1 vccd1 _16005_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_94_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1172 _15946_/A2 vssd1 vssd1 vccd1 vccd1 _15910_/A2 sky130_fd_sc_hd__buf_4
X_17846_ _19319_/CLK _17846_/D vssd1 vssd1 vccd1 vccd1 _17846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1183 _15526_/B vssd1 vssd1 vccd1 vccd1 _15404_/B sky130_fd_sc_hd__buf_4
XFILLER_282_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1194 _16969_/B1 vssd1 vssd1 vccd1 vccd1 _16965_/B1 sky130_fd_sc_hd__buf_4
XFILLER_67_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14989_ _15009_/A1 _18272_/Q _14988_/Y _11712_/A vssd1 vssd1 vccd1 vccd1 _14989_/X
+ sky130_fd_sc_hd__a31o_1
X_17777_ _19573_/CLK _17777_/D vssd1 vssd1 vccd1 vccd1 _17777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19516_ _19521_/CLK _19516_/D vssd1 vssd1 vccd1 vccd1 _19516_/Q sky130_fd_sc_hd__dfxtp_1
X_16728_ _19262_/Q _19261_/Q _16728_/C vssd1 vssd1 vccd1 vccd1 _16734_/C sky130_fd_sc_hd__and3_1
XFILLER_34_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16659_ _16768_/A _16659_/B _16664_/C vssd1 vssd1 vccd1 vccd1 _19241_/D sky130_fd_sc_hd__nor3_1
XFILLER_222_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19447_ _19482_/CLK _19447_/D vssd1 vssd1 vccd1 vccd1 _19447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09200_ _10282_/A1 _18143_/Q _18789_/Q _10141_/S _10293_/B1 vssd1 vssd1 vccd1 vccd1
+ _09200_/X sky130_fd_sc_hd__a221o_1
XFILLER_167_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19378_ _19540_/CLK _19378_/D vssd1 vssd1 vccd1 vccd1 _19378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09131_ _19078_/Q _18982_/Q _09269_/S vssd1 vssd1 vccd1 vccd1 _09131_/X sky130_fd_sc_hd__mux2_1
X_18329_ _19211_/CLK _18329_/D vssd1 vssd1 vccd1 vccd1 _18329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09062_ _17892_/Q _09062_/B _17893_/Q vssd1 vssd1 vccd1 vccd1 _12261_/B sky130_fd_sc_hd__and3b_1
XFILLER_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_96_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19140_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_25_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19197_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_265_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09964_ _10747_/A1 _09963_/X _08903_/A vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__a21o_1
XFILLER_170_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08915_ _08816_/A _16392_/B vssd1 vssd1 vccd1 vccd1 _14350_/A sky130_fd_sc_hd__nand2b_4
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09895_ _09367_/B _15130_/A _09866_/Y vssd1 vssd1 vccd1 vccd1 _12602_/B sky130_fd_sc_hd__a21bo_4
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08846_ _09708_/A vssd1 vssd1 vccd1 vccd1 _08846_/Y sky130_fd_sc_hd__inv_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_506 _14423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_517 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_528 _11719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_539 input238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10670_ _10589_/S _10665_/Y _10669_/Y _11602_/C1 vssd1 vssd1 vccd1 vccd1 _10670_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ input169/X input141/X _09990_/S vssd1 vssd1 vccd1 vccd1 _09329_/X sky130_fd_sc_hd__mux2_8
XFILLER_167_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12340_ _12382_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _12340_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12271_ _12271_/A _12271_/B vssd1 vssd1 vccd1 vccd1 _12277_/A sky130_fd_sc_hd__or2_1
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14010_ _17970_/Q _14028_/A vssd1 vssd1 vccd1 vccd1 _14010_/X sky130_fd_sc_hd__or2_1
XFILLER_181_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11222_ _09987_/A _11221_/X _11216_/X vssd1 vssd1 vccd1 vccd1 _11222_/X sky130_fd_sc_hd__o21a_1
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11153_ _18423_/Q _11224_/B _11152_/X _10706_/S vssd1 vssd1 vccd1 vccd1 _11153_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10104_ _18163_/Q _11482_/A2 _10103_/X _11406_/B2 vssd1 vssd1 vccd1 vccd1 _10104_/X
+ sky130_fd_sc_hd__a211o_1
X_15961_ _18696_/Q _15977_/A2 _15960_/X _16892_/A vssd1 vssd1 vccd1 vccd1 _18696_/D
+ sky130_fd_sc_hd__o211a_1
X_11084_ _11082_/X _11083_/X _11084_/S vssd1 vssd1 vccd1 vccd1 _11084_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput220 localMemory_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input220/X sky130_fd_sc_hd__clkbuf_16
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput231 localMemory_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 input231/X sky130_fd_sc_hd__buf_12
XFILLER_249_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17700_ _17700_/A0 _19626_/Q _17722_/S vssd1 vssd1 vccd1 vccd1 _19626_/D sky130_fd_sc_hd__mux2_1
Xinput242 localMemory_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input242/X sky130_fd_sc_hd__buf_8
X_14912_ _14912_/A1 _13659_/X _14983_/B1 _18648_/Q _14973_/C1 vssd1 vssd1 vccd1 vccd1
+ _14912_/X sky130_fd_sc_hd__a221o_1
X_10035_ _11618_/A1 _18133_/Q _18779_/Q _11609_/S vssd1 vssd1 vccd1 vccd1 _10035_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput253 manufacturerID[0] vssd1 vssd1 vccd1 vccd1 _15857_/A sky130_fd_sc_hd__buf_4
X_18680_ _18683_/CLK _18680_/D vssd1 vssd1 vccd1 vccd1 _18680_/Q sky130_fd_sc_hd__dfxtp_1
X_15892_ _18673_/Q _15910_/A2 _15891_/X _15904_/C1 vssd1 vssd1 vccd1 vccd1 _18673_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_236_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput264 partID[0] vssd1 vssd1 vccd1 vccd1 _15890_/A sky130_fd_sc_hd__buf_2
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput275 partID[5] vssd1 vssd1 vccd1 vccd1 _15905_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_264_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ _17664_/A0 _19559_/Q _17654_/S vssd1 vssd1 vccd1 vccd1 _19559_/D sky130_fd_sc_hd__mux2_1
X_14843_ _14865_/A1 _14842_/X _14865_/B1 vssd1 vssd1 vccd1 vccd1 _14843_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_48_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17562_ _17123_/B _17583_/B _17588_/B1 _17561_/X vssd1 vssd1 vccd1 vccd1 _19523_/D
+ sky130_fd_sc_hd__o211a_1
X_14774_ input105/X input77/X _14784_/S vssd1 vssd1 vccd1 vccd1 _14775_/A sky130_fd_sc_hd__mux2_1
XFILLER_251_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11986_ _14074_/B _16459_/B vssd1 vssd1 vccd1 vccd1 _14272_/B sky130_fd_sc_hd__or2_4
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19301_ _19326_/CLK _19301_/D vssd1 vssd1 vccd1 vccd1 _19301_/Q sky130_fd_sc_hd__dfxtp_1
X_16513_ _17679_/A0 _19119_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _19119_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13725_ _13930_/A1 _13711_/Y _13930_/B1 vssd1 vssd1 vccd1 vccd1 _13725_/X sky130_fd_sc_hd__o21a_1
X_17493_ _17493_/A _17493_/B vssd1 vssd1 vccd1 vccd1 _17493_/Y sky130_fd_sc_hd__nand2_1
X_10937_ _18255_/Q _10940_/S _10633_/A _10936_/X vssd1 vssd1 vccd1 vccd1 _10937_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19232_ _19268_/CLK _19232_/D vssd1 vssd1 vccd1 vccd1 _19232_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16444_ _19052_/Q _16609_/A0 _16453_/S vssd1 vssd1 vccd1 vccd1 _19052_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13656_ _19350_/Q _13950_/A2 _13950_/B1 _19478_/Q _13950_/C1 vssd1 vssd1 vccd1 vccd1
+ _13656_/X sky130_fd_sc_hd__a221o_1
X_10868_ _10841_/X _10844_/X _10399_/A vssd1 vssd1 vccd1 vccd1 _10868_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12607_ _12957_/A _12957_/B _12601_/Y vssd1 vssd1 vccd1 vccd1 _12985_/B sky130_fd_sc_hd__o21a_1
X_19163_ _19163_/CLK _19163_/D vssd1 vssd1 vccd1 vccd1 _19163_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _17674_/A0 _18986_/Q _16385_/S vssd1 vssd1 vccd1 vccd1 _18986_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _19510_/Q _13947_/A2 _13947_/B1 _13586_/X vssd1 vssd1 vccd1 vccd1 _13587_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10799_ _18037_/Q _18005_/Q _11604_/S vssd1 vssd1 vccd1 vccd1 _10799_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18114_ _19450_/CLK _18114_/D vssd1 vssd1 vccd1 vccd1 _18114_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_157_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ _17129_/A _15325_/X _15424_/C1 vssd1 vssd1 vccd1 vccd1 _15326_/X sky130_fd_sc_hd__a21o_1
X_19094_ _19596_/CLK _19094_/D vssd1 vssd1 vccd1 vccd1 _19094_/Q sky130_fd_sc_hd__dfxtp_1
X_12538_ _12538_/A _12538_/B vssd1 vssd1 vccd1 vccd1 _12538_/Y sky130_fd_sc_hd__nor2_2
XFILLER_129_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18045_ _19615_/CLK _18045_/D vssd1 vssd1 vccd1 vccd1 _18045_/Q sky130_fd_sc_hd__dfxtp_1
X_15257_ _18569_/Q _15351_/A2 _15251_/X _15256_/X _17338_/A vssd1 vssd1 vccd1 vccd1
+ _18569_/D sky130_fd_sc_hd__o221a_1
X_12469_ _16852_/A _14675_/C _12468_/Y vssd1 vssd1 vccd1 vccd1 _12851_/B sky130_fd_sc_hd__o21a_4
X_14208_ _18102_/Q _14266_/B vssd1 vssd1 vccd1 vccd1 _14208_/X sky130_fd_sc_hd__or2_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15188_ _15186_/Y _15188_/B vssd1 vssd1 vccd1 vccd1 _15189_/B sky130_fd_sc_hd__and2b_1
XFILLER_259_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14139_ _15832_/A1 _18078_/Q _14139_/S vssd1 vssd1 vccd1 vccd1 _18078_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18947_ _19564_/CLK _18947_/D vssd1 vssd1 vccd1 vccd1 _18947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09680_ _12468_/B _18208_/Q _09680_/B1 _18943_/Q vssd1 vssd1 vccd1 vccd1 _09680_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18878_ _19589_/CLK _18878_/D vssd1 vssd1 vccd1 vccd1 _18878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_143_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17814_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_282_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17829_ _19306_/CLK _17829_/D vssd1 vssd1 vccd1 vccd1 _17829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09114_ _18418_/Q _11479_/B _09129_/S _09113_/X vssd1 vssd1 vccd1 vccd1 _09114_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09045_ _09652_/A _09045_/B vssd1 vssd1 vccd1 vccd1 _09046_/B sky130_fd_sc_hd__nor2_1
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1908 _11712_/A vssd1 vssd1 vccd1 vccd1 _14928_/B1 sky130_fd_sc_hd__clkbuf_2
Xfanout910 _16425_/S vssd1 vssd1 vccd1 vccd1 _16421_/S sky130_fd_sc_hd__buf_12
XFILLER_278_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout921 _16255_/S vssd1 vssd1 vccd1 vccd1 _16258_/S sky130_fd_sc_hd__clkbuf_16
X_09947_ _12933_/A vssd1 vssd1 vccd1 vccd1 _09947_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout932 _15083_/Y vssd1 vssd1 vccd1 vccd1 _17445_/B1 sky130_fd_sc_hd__buf_2
Xfanout943 _14994_/B vssd1 vssd1 vccd1 vccd1 _14893_/S sky130_fd_sc_hd__buf_4
Xfanout954 _14599_/X vssd1 vssd1 vccd1 vccd1 _14622_/S sky130_fd_sc_hd__buf_4
XFILLER_277_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout965 _14075_/Y vssd1 vssd1 vccd1 vccd1 _14107_/S sky130_fd_sc_hd__buf_12
Xfanout976 _13527_/B1 vssd1 vssd1 vccd1 vccd1 _13920_/B2 sky130_fd_sc_hd__buf_4
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout987 _13973_/A2 vssd1 vssd1 vccd1 vccd1 _13940_/A2 sky130_fd_sc_hd__buf_2
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _18309_/Q _17760_/Q _09885_/S vssd1 vssd1 vccd1 vccd1 _09878_/X sky130_fd_sc_hd__mux2_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout998 _17684_/A0 vssd1 vssd1 vccd1 vccd1 _16551_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_245_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08829_ _18590_/Q vssd1 vssd1 vccd1 vccd1 _17533_/A sky130_fd_sc_hd__inv_2
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 _18112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11840_ _11844_/A _11840_/B vssd1 vssd1 vccd1 vccd1 _11840_/X sky130_fd_sc_hd__and2_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_314 _18102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_325 _18109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_336 wire989/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_347 fanout1525/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_358 _12461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11771_ _13810_/A _11730_/Y _14522_/A2 _18589_/Q vssd1 vssd1 vccd1 vccd1 _11771_/X
+ sky130_fd_sc_hd__a2bb2o_4
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_369 _14487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ _13970_/B2 _13482_/A _13509_/X _13899_/A vssd1 vssd1 vccd1 vccd1 _13511_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10722_ _18648_/Q _10726_/S vssd1 vssd1 vccd1 vccd1 _10722_/X sky130_fd_sc_hd__or2_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _17692_/A0 _18340_/Q _14521_/S vssd1 vssd1 vccd1 vccd1 _18340_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13441_ _13936_/B2 _13408_/A _13440_/X _15429_/A2 vssd1 vssd1 vccd1 vccd1 _13442_/B
+ sky130_fd_sc_hd__a22o_1
X_10653_ _10653_/A1 _10645_/X _10644_/X _10653_/C1 vssd1 vssd1 vccd1 vccd1 _10653_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_22_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16160_ _18276_/D _16156_/B _16159_/X vssd1 vssd1 vccd1 vccd1 _18778_/D sky130_fd_sc_hd__a21o_1
XFILLER_166_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13372_ _19536_/Q _19504_/Q _13372_/S vssd1 vssd1 vccd1 vccd1 _13372_/X sky130_fd_sc_hd__mux2_1
X_10584_ _10662_/A1 _19219_/Q _19187_/Q _10645_/S _08899_/A vssd1 vssd1 vccd1 vccd1
+ _10584_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15111_ _15111_/A _15133_/B vssd1 vssd1 vccd1 vccd1 _15112_/B sky130_fd_sc_hd__nand2_4
X_12323_ _12323_/A _12323_/B vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__or2_4
X_16091_ _18748_/Q _16093_/B vssd1 vssd1 vccd1 vccd1 _16091_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15042_ _18530_/Q _14666_/X _18531_/Q vssd1 vssd1 vccd1 vccd1 _15043_/C sky130_fd_sc_hd__o21ai_1
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12254_ _16808_/A _12256_/B vssd1 vssd1 vccd1 vccd1 _12254_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11205_ _11203_/X _11204_/X _11285_/S vssd1 vssd1 vccd1 vccd1 _11205_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12185_ _12187_/A _12185_/B _12186_/B vssd1 vssd1 vccd1 vccd1 _17858_/D sky130_fd_sc_hd__nor3_1
XFILLER_123_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18801_ _19025_/CLK _18801_/D vssd1 vssd1 vccd1 vccd1 _18801_/Q sky130_fd_sc_hd__dfxtp_1
X_11136_ _11138_/B vssd1 vssd1 vccd1 vccd1 _11136_/Y sky130_fd_sc_hd__clkinv_2
X_16993_ _19333_/Q _17043_/B vssd1 vssd1 vccd1 vccd1 _16993_/X sky130_fd_sc_hd__or2_1
XFILLER_283_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18732_ _18734_/CLK _18732_/D vssd1 vssd1 vccd1 vccd1 _18732_/Q sky130_fd_sc_hd__dfxtp_1
X_15944_ input7/X _12851_/A _15947_/S vssd1 vssd1 vccd1 vccd1 _15944_/X sky130_fd_sc_hd__mux2_1
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11067_ _17937_/Q _11451_/A2 _11066_/Y _08947_/B vssd1 vssd1 vccd1 vccd1 _11067_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_95_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10018_ _11566_/A1 _19195_/Q _19163_/Q _11226_/S _09086_/A vssd1 vssd1 vccd1 vccd1
+ _10020_/B sky130_fd_sc_hd__a221o_1
X_18663_ _18666_/CLK _18663_/D vssd1 vssd1 vccd1 vccd1 _18663_/Q sky130_fd_sc_hd__dfxtp_1
X_15875_ _15875_/A _15905_/B _15908_/C vssd1 vssd1 vccd1 vccd1 _15875_/X sky130_fd_sc_hd__and3_1
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _15009_/A1 _18270_/Q _14825_/Y _14918_/B1 vssd1 vssd1 vccd1 vccd1 _14826_/X
+ sky130_fd_sc_hd__a31o_2
X_17614_ _19548_/Q _17624_/A2 _17613_/X _17592_/B vssd1 vssd1 vccd1 vccd1 _19548_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18594_ _18875_/CLK _18594_/D vssd1 vssd1 vccd1 vccd1 _18594_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ _14754_/Y _14756_/Y _14879_/B1 vssd1 vssd1 vccd1 vccd1 _14757_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17545_ _18592_/Q _17550_/A _17544_/X _17545_/C1 vssd1 vssd1 vccd1 vccd1 _17545_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_251_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11969_ _18739_/Q _16034_/S vssd1 vssd1 vccd1 vccd1 _16041_/A sky130_fd_sc_hd__nand2_4
XFILLER_204_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13708_ _13739_/A _13695_/A _13707_/X vssd1 vssd1 vccd1 vccd1 _13708_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_260_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17476_ _18579_/Q _17527_/A1 _17516_/C1 vssd1 vssd1 vccd1 vccd1 _17476_/X sky130_fd_sc_hd__o21a_1
XFILLER_189_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14688_ _14688_/A _14688_/B _14688_/C _14688_/D vssd1 vssd1 vccd1 vccd1 _15834_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_204_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19215_ _19575_/CLK _19215_/D vssd1 vssd1 vccd1 vccd1 _19215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13639_ _13638_/B _13637_/X _13638_/Y _13930_/B1 _13931_/A vssd1 vssd1 vccd1 vccd1
+ _13639_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16427_ _19035_/Q _17692_/A0 _16458_/S vssd1 vssd1 vccd1 vccd1 _19035_/D sky130_fd_sc_hd__mux2_1
XFILLER_220_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16358_ _18970_/Q _16557_/A0 _16358_/S vssd1 vssd1 vccd1 vccd1 _18970_/D sky130_fd_sc_hd__mux2_1
X_19146_ _19146_/CLK _19146_/D vssd1 vssd1 vccd1 vccd1 _19146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15309_ _15289_/A _15289_/B _15293_/B vssd1 vssd1 vccd1 vccd1 _15310_/B sky130_fd_sc_hd__a21o_1
X_19077_ _19564_/CLK _19077_/D vssd1 vssd1 vccd1 vccd1 _19077_/Q sky130_fd_sc_hd__dfxtp_1
X_16289_ _16455_/A1 _18903_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _18903_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18028_ _19630_/CLK _18028_/D vssd1 vssd1 vccd1 vccd1 _18028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09801_ _18019_/Q _17987_/Q _09801_/S vssd1 vssd1 vccd1 vccd1 _09801_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09732_ _14214_/A _15173_/A _09948_/B vssd1 vssd1 vccd1 vccd1 _12609_/B sky130_fd_sc_hd__mux2_8
XFILLER_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09663_ _18847_/Q _18879_/Q _09671_/S vssd1 vssd1 vccd1 vccd1 _09663_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09594_ _18537_/Q _18412_/Q _10362_/S vssd1 vssd1 vccd1 vccd1 _09594_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19211_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09028_ _09043_/A _09028_/B vssd1 vssd1 vccd1 vccd1 _09986_/B sky130_fd_sc_hd__nor2_2
XFILLER_3_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1705 _08843_/Y vssd1 vssd1 vccd1 vccd1 _09086_/A sky130_fd_sc_hd__buf_12
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1716 _16898_/A1 vssd1 vssd1 vccd1 vccd1 _12492_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_160_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1727 _16969_/C1 vssd1 vssd1 vccd1 vccd1 _16965_/C1 sky130_fd_sc_hd__buf_4
XFILLER_265_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1738 _15009_/A1 vssd1 vssd1 vccd1 vccd1 _14696_/A sky130_fd_sc_hd__buf_6
Xfanout740 _16607_/A0 vssd1 vssd1 vccd1 vccd1 _17707_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_278_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1749 _17921_/Q vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__buf_6
Xfanout751 _09816_/A vssd1 vssd1 vccd1 vccd1 _13046_/A1 sky130_fd_sc_hd__buf_4
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout762 _16471_/A0 vssd1 vssd1 vccd1 vccd1 _17670_/A0 sky130_fd_sc_hd__clkbuf_4
X_13990_ _14032_/B _13990_/B vssd1 vssd1 vccd1 vccd1 _13990_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout773 _17625_/Y vssd1 vssd1 vccd1 vccd1 _17657_/S sky130_fd_sc_hd__buf_12
XFILLER_283_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout784 _16558_/Y vssd1 vssd1 vccd1 vccd1 _16590_/S sky130_fd_sc_hd__buf_8
Xfanout795 _16355_/S vssd1 vssd1 vccd1 vccd1 _16357_/S sky130_fd_sc_hd__buf_12
XFILLER_74_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _13129_/B _13130_/B _13089_/A vssd1 vssd1 vccd1 vccd1 _12941_/X sky130_fd_sc_hd__mux2_2
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _15744_/A _15687_/A _15645_/B vssd1 vssd1 vccd1 vccd1 _15665_/B sky130_fd_sc_hd__a21o_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _12942_/S _12872_/B vssd1 vssd1 vccd1 vccd1 _12872_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_100 _11067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _11751_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _17670_/A0 _18418_/Q _14630_/S vssd1 vssd1 vccd1 vccd1 _18418_/D sky130_fd_sc_hd__mux2_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_122 _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_133 _11814_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ _11823_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11858_/B sky130_fd_sc_hd__nor2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15591_/A _15591_/B vssd1 vssd1 vccd1 vccd1 _15591_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_60_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_144 _11868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _11872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_166 _13024_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17330_ _17330_/A _17330_/B vssd1 vssd1 vccd1 vccd1 _19462_/D sky130_fd_sc_hd__nor2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _14002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ _14596_/A _14542_/B vssd1 vssd1 vccd1 vccd1 _18379_/D sky130_fd_sc_hd__or2_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_188 _13709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _18572_/Q _11726_/B _11799_/B _13224_/A vssd1 vssd1 vccd1 vccd1 _11754_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_199 _13939_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17261_ _17261_/A _17261_/B vssd1 vssd1 vccd1 vccd1 _19437_/D sky130_fd_sc_hd__nor2_1
X_10705_ _11250_/A1 _19153_/Q _11154_/S _19121_/Q vssd1 vssd1 vccd1 vccd1 _10705_/X
+ sky130_fd_sc_hd__o22a_1
X_14473_ _18325_/Q _17677_/A0 _14485_/S vssd1 vssd1 vccd1 vccd1 _18325_/D sky130_fd_sc_hd__mux2_1
X_11685_ _13566_/A _13545_/B _13512_/B _11685_/D vssd1 vssd1 vccd1 vccd1 _11686_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_202_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19000_ _19613_/CLK _19000_/D vssd1 vssd1 vccd1 vccd1 _19000_/Q sky130_fd_sc_hd__dfxtp_1
X_16212_ _17709_/A0 _18828_/Q _16212_/S vssd1 vssd1 vccd1 vccd1 _18828_/D sky130_fd_sc_hd__mux2_1
X_13424_ _17838_/Q _13821_/B _12548_/X vssd1 vssd1 vccd1 vccd1 _13424_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17192_ _17198_/A _17192_/B vssd1 vssd1 vccd1 vccd1 _19415_/D sky130_fd_sc_hd__nor2_1
X_10636_ _10633_/X _10635_/X _10629_/X vssd1 vssd1 vccd1 vccd1 _10636_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_220_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16143_ _18776_/Q _16143_/B _16143_/C _18775_/Q vssd1 vssd1 vccd1 vccd1 _16154_/A
+ sky130_fd_sc_hd__or4b_2
X_13355_ _13354_/A _13038_/B _13354_/Y _13194_/S vssd1 vssd1 vccd1 vccd1 _13355_/X
+ sky130_fd_sc_hd__o211a_1
X_10567_ _18556_/Q _18431_/Q _10645_/S vssd1 vssd1 vccd1 vccd1 _10567_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ _16852_/A _14687_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _16819_/B sky130_fd_sc_hd__or3b_4
X_16074_ _18741_/Q _11981_/B _16063_/C _16075_/A vssd1 vssd1 vccd1 vccd1 _16074_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13286_ _13928_/A1 _13275_/X _13285_/X vssd1 vssd1 vccd1 vccd1 _13996_/B sky130_fd_sc_hd__a21oi_4
XFILLER_154_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10498_ _19124_/Q _19156_/Q _10500_/S vssd1 vssd1 vccd1 vccd1 _10498_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15025_ _18514_/Q input191/X _15038_/S vssd1 vssd1 vccd1 vccd1 _18514_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ _17878_/Q _12240_/C _12241_/A vssd1 vssd1 vccd1 vccd1 _12237_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_142_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12168_ _17851_/Q _17852_/Q _12168_/C vssd1 vssd1 vccd1 vccd1 _12170_/B sky130_fd_sc_hd__and3_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11119_ _11352_/A1 _18150_/Q _18796_/Q _11125_/B2 vssd1 vssd1 vccd1 vccd1 _11119_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_283_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12099_ _17826_/Q _12100_/C _12098_/Y vssd1 vssd1 vccd1 vccd1 _17826_/D sky130_fd_sc_hd__o21a_1
X_16976_ _17047_/B vssd1 vssd1 vccd1 vccd1 _16977_/B sky130_fd_sc_hd__clkinv_2
XFILLER_284_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18715_ _18715_/CLK _18715_/D vssd1 vssd1 vccd1 vccd1 _18715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 coreIndex[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_6
X_15927_ _18684_/Q _15948_/A2 _15923_/C _15926_/X _15945_/C1 vssd1 vssd1 vccd1 vccd1
+ _15927_/X sky130_fd_sc_hd__a221o_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18646_ _19611_/CLK _18646_/D vssd1 vssd1 vccd1 vccd1 _18646_/Q sky130_fd_sc_hd__dfxtp_4
X_15858_ _18661_/Q _15853_/Y _15906_/B1 vssd1 vssd1 vccd1 vccd1 _15858_/X sky130_fd_sc_hd__a21o_1
XFILLER_252_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14809_ _12459_/X _13998_/B _14683_/X _18638_/Q vssd1 vssd1 vccd1 vccd1 _14809_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18577_ _19531_/CLK _18577_/D vssd1 vssd1 vccd1 vccd1 _18577_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_224_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15789_ _15789_/A1 _15788_/Y _15789_/B1 vssd1 vssd1 vccd1 vccd1 _15789_/X sky130_fd_sc_hd__a21o_1
XFILLER_205_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17528_ _18128_/Q _17528_/B vssd1 vssd1 vccd1 vccd1 _17528_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17459_ _19503_/Q _17462_/B _17458_/X _17338_/A vssd1 vssd1 vccd1 vccd1 _19503_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_193_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19129_ _19628_/CLK _19129_/D vssd1 vssd1 vccd1 vccd1 _19129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput310 _11758_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[14] sky130_fd_sc_hd__buf_4
XFILLER_105_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput321 _11768_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[24] sky130_fd_sc_hd__buf_4
XFILLER_160_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput332 _11752_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[9] sky130_fd_sc_hd__buf_4
XFILLER_160_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput343 _11849_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[18] sky130_fd_sc_hd__buf_4
Xoutput354 _11894_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[28] sky130_fd_sc_hd__buf_4
XFILLER_236_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput365 _11810_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[9] sky130_fd_sc_hd__buf_4
Xoutput376 _11920_/X vssd1 vssd1 vccd1 vccd1 din0[0] sky130_fd_sc_hd__buf_4
XFILLER_0_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput387 _11921_/X vssd1 vssd1 vccd1 vccd1 din0[1] sky130_fd_sc_hd__buf_4
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput398 _11922_/X vssd1 vssd1 vccd1 vccd1 din0[2] sky130_fd_sc_hd__buf_4
XFILLER_248_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09715_ _10747_/A1 _09714_/X _09709_/X _08903_/A vssd1 vssd1 vccd1 vccd1 _09715_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_228_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09646_ _12614_/B _09647_/B vssd1 vssd1 vccd1 vccd1 _09648_/B sky130_fd_sc_hd__nor2_1
XFILLER_255_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _10366_/A1 _19200_/Q _19168_/Q _10362_/S _12766_/A0 vssd1 vssd1 vccd1 vccd1
+ _09577_/X sky130_fd_sc_hd__a221o_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ _11478_/S _11470_/B vssd1 vssd1 vccd1 vccd1 _11470_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10421_ _18042_/Q _18010_/Q _10424_/S vssd1 vssd1 vccd1 vccd1 _10421_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13140_ _13194_/S _13139_/Y _13197_/B1 vssd1 vssd1 vccd1 vccd1 _13140_/X sky130_fd_sc_hd__a21o_1
X_10352_ _10205_/S _10351_/X _10350_/X _11046_/S1 vssd1 vssd1 vccd1 vccd1 _10352_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ input7/X _12552_/X _13070_/X _12538_/B vssd1 vssd1 vccd1 vccd1 _13071_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_140_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10283_ _10275_/S _10281_/X _10282_/X _09429_/S vssd1 vssd1 vccd1 vccd1 _10283_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12022_ _17789_/Q _17690_/A0 _12022_/S vssd1 vssd1 vccd1 vccd1 _17789_/D sky130_fd_sc_hd__mux2_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1502 _08968_/S0 vssd1 vssd1 vccd1 vccd1 _09498_/S sky130_fd_sc_hd__clkbuf_4
Xfanout1513 fanout1514/X vssd1 vssd1 vccd1 vccd1 _10199_/S sky130_fd_sc_hd__buf_4
XFILLER_160_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1524 fanout1525/X vssd1 vssd1 vccd1 vccd1 fanout1524/X sky130_fd_sc_hd__buf_4
XFILLER_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16830_ _16821_/A _17818_/Q _12474_/Y vssd1 vssd1 vccd1 vccd1 _16831_/B sky130_fd_sc_hd__a21o_1
Xfanout1535 _10653_/A1 vssd1 vssd1 vccd1 vccd1 _09976_/A1 sky130_fd_sc_hd__buf_4
XFILLER_265_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1546 _11616_/S vssd1 vssd1 vccd1 vccd1 _10040_/S sky130_fd_sc_hd__buf_6
XFILLER_116_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1557 _09381_/S vssd1 vssd1 vccd1 vccd1 _11428_/A sky130_fd_sc_hd__buf_6
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1568 _11495_/B1 vssd1 vssd1 vccd1 vccd1 _11417_/B1 sky130_fd_sc_hd__buf_12
XFILLER_219_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout570 _15124_/C vssd1 vssd1 vccd1 vccd1 _15133_/B sky130_fd_sc_hd__buf_8
XFILLER_93_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1579 fanout1581/X vssd1 vssd1 vccd1 vccd1 _11507_/S sky130_fd_sc_hd__buf_8
Xfanout581 _12412_/A vssd1 vssd1 vccd1 vccd1 _12430_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout592 _14247_/A2 vssd1 vssd1 vccd1 vccd1 _14267_/A2 sky130_fd_sc_hd__buf_4
XFILLER_93_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16761_ _19274_/Q _16762_/B vssd1 vssd1 vccd1 vccd1 _16763_/B sky130_fd_sc_hd__nor2_1
XFILLER_247_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13973_ _17951_/Q _13973_/A2 _13971_/X _13972_/Y _15039_/A vssd1 vssd1 vccd1 vccd1
+ _17951_/D sky130_fd_sc_hd__o221a_1
XFILLER_281_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18500_ _18501_/CLK _18500_/D vssd1 vssd1 vccd1 vccd1 _18500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15712_ _19483_/Q _19417_/Q vssd1 vssd1 vccd1 vccd1 _15713_/B sky130_fd_sc_hd__nand2_1
X_12924_ _13438_/A _12906_/X _13956_/B1 vssd1 vssd1 vccd1 vccd1 _12924_/X sky130_fd_sc_hd__a21o_1
X_16692_ _19250_/Q _16695_/C _12203_/A vssd1 vssd1 vccd1 vccd1 _16692_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_234_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19480_ _19483_/CLK _19480_/D vssd1 vssd1 vccd1 vccd1 _19480_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_234_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18431_ _19638_/CLK _18431_/D vssd1 vssd1 vccd1 vccd1 _18431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12855_ _19330_/Q _12578_/Y _12853_/X _12854_/X _12529_/Y vssd1 vssd1 vccd1 vccd1
+ _12855_/X sky130_fd_sc_hd__a221o_1
X_15643_ _15686_/A _15644_/B vssd1 vssd1 vccd1 vccd1 _15645_/A sky130_fd_sc_hd__and2_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11806_ _11810_/A _11818_/B _11806_/C vssd1 vssd1 vccd1 vccd1 _11806_/X sky130_fd_sc_hd__and3_1
X_18362_ _19025_/CLK _18362_/D vssd1 vssd1 vccd1 vccd1 _18362_/Q sky130_fd_sc_hd__dfxtp_1
X_15574_ _13643_/X _15110_/X _10828_/Y _15111_/A vssd1 vssd1 vccd1 vccd1 _15574_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12786_ _17889_/Q _17888_/Q _15082_/A vssd1 vssd1 vccd1 vccd1 _12786_/X sky130_fd_sc_hd__a21o_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _19455_/Q _17313_/B vssd1 vssd1 vccd1 vccd1 _17313_/Y sky130_fd_sc_hd__nand2_1
X_14525_ _14525_/A _14525_/B _14596_/A vssd1 vssd1 vccd1 vccd1 _18372_/D sky130_fd_sc_hd__nor3_1
XFILLER_109_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _12985_/A _11737_/B vssd1 vssd1 vccd1 vccd1 _11737_/X sky130_fd_sc_hd__xor2_4
XFILLER_175_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18293_ _18593_/CLK _18293_/D vssd1 vssd1 vccd1 vccd1 _18293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14456_ _18308_/Q _17660_/A0 _14483_/S vssd1 vssd1 vccd1 vccd1 _18308_/D sky130_fd_sc_hd__mux2_1
X_17244_ _19432_/Q _17244_/B vssd1 vssd1 vccd1 vccd1 _17244_/Y sky130_fd_sc_hd__nand2_1
X_11668_ _13695_/A vssd1 vssd1 vccd1 vccd1 _11668_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13407_ _13479_/C _13407_/B vssd1 vssd1 vccd1 vccd1 _13408_/A sky130_fd_sc_hd__or2_1
XFILLER_179_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10619_ _18866_/Q _18898_/Q _10619_/S vssd1 vssd1 vccd1 vccd1 _10619_/X sky130_fd_sc_hd__mux2_1
X_17175_ _17214_/A _17175_/B vssd1 vssd1 vccd1 vccd1 _17483_/A sky130_fd_sc_hd__nand2_1
X_14387_ _17661_/A0 _18238_/Q _14402_/S vssd1 vssd1 vccd1 vccd1 _18238_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11599_ _11597_/X _11598_/X _11606_/S vssd1 vssd1 vccd1 vccd1 _11599_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16126_ _16140_/A1 _16125_/Y _16128_/B1 vssd1 vssd1 vccd1 vccd1 _18765_/D sky130_fd_sc_hd__a21oi_1
XFILLER_115_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13338_ _19437_/Q _12582_/X _13337_/X vssd1 vssd1 vccd1 vccd1 _13338_/X sky130_fd_sc_hd__o21a_2
XFILLER_127_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16057_ _16063_/A _16055_/A _16041_/X _14164_/B vssd1 vssd1 vccd1 vccd1 _16057_/X
+ sky130_fd_sc_hd__o211a_1
X_13269_ _14154_/B1 _13266_/X _13268_/X _09145_/A _13262_/X vssd1 vssd1 vccd1 vccd1
+ _13269_/X sky130_fd_sc_hd__o221a_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ _15008_/A vssd1 vssd1 vccd1 vccd1 _15008_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16959_ _19324_/Q _17205_/B _16963_/S vssd1 vssd1 vccd1 vccd1 _16960_/B sky130_fd_sc_hd__mux2_1
XFILLER_271_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09500_ _09495_/X _09496_/X _10301_/S vssd1 vssd1 vccd1 vccd1 _09500_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09431_ _09426_/Y _09430_/Y _11516_/B1 vssd1 vssd1 vccd1 vccd1 _09431_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18629_ _19211_/CLK _18629_/D vssd1 vssd1 vccd1 vccd1 _18629_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09362_ _11459_/B1 _09347_/X _09360_/X _09361_/X vssd1 vssd1 vccd1 vccd1 _09362_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09293_ _18448_/Q _18349_/Q _09302_/S vssd1 vssd1 vccd1 vccd1 _09293_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_11 _14718_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_22 _14990_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 _08899_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_44 _12600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_55 _09743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_66 _13874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_77 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_88 _10459_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_99 _11067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10970_ _18551_/Q _18426_/Q _18035_/Q _18003_/Q _11340_/B2 _11357_/S1 vssd1 vssd1
+ vccd1 vccd1 _10970_/X sky130_fd_sc_hd__mux4_1
XFILLER_216_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09629_ _09627_/X _09628_/X _11161_/S vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__mux2_1
XFILLER_189_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _10832_/A _12640_/B vssd1 vssd1 vccd1 vccd1 _12640_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_62_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12571_ _13246_/B1 _13243_/B1 _12570_/X _12568_/Y vssd1 vssd1 vccd1 vccd1 _12571_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _18167_/Q _17694_/A0 _14339_/S vssd1 vssd1 vccd1 vccd1 _18167_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11522_ _12625_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11523_/B sky130_fd_sc_hd__nor2_2
XFILLER_196_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15290_ _15290_/A _15310_/A vssd1 vssd1 vccd1 vccd1 _15365_/B sky130_fd_sc_hd__and2_1
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14241_ _18292_/Q _14267_/A2 _14240_/X _14452_/B vssd1 vssd1 vccd1 vccd1 _18118_/D
+ sky130_fd_sc_hd__o211a_1
X_11453_ _18983_/Q _11479_/B vssd1 vssd1 vccd1 vccd1 _11453_/X sky130_fd_sc_hd__or2_1
XFILLER_137_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ _09129_/S _10403_/X _11466_/B1 vssd1 vssd1 vccd1 vccd1 _10404_/X sky130_fd_sc_hd__o21a_1
X_14172_ _18697_/Q _18084_/Q _14186_/S vssd1 vssd1 vccd1 vccd1 _14173_/B sky130_fd_sc_hd__mux2_1
X_11384_ _18545_/Q _11384_/B vssd1 vssd1 vccd1 vccd1 _11384_/X sky130_fd_sc_hd__or2_1
XFILLER_124_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13123_ _13079_/A _13119_/Y _13120_/X _13125_/A _13254_/B2 vssd1 vssd1 vccd1 vccd1
+ _13123_/X sky130_fd_sc_hd__a32o_1
X_10335_ _10333_/X _10334_/X _10335_/S vssd1 vssd1 vccd1 vccd1 _10336_/B sky130_fd_sc_hd__mux2_1
XFILLER_180_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18980_ _19076_/CLK _18980_/D vssd1 vssd1 vccd1 vccd1 _18980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _17931_/CLK _17931_/D vssd1 vssd1 vccd1 vccd1 _17931_/Q sky130_fd_sc_hd__dfxtp_4
X_13054_ _18107_/Q _13055_/B vssd1 vssd1 vccd1 vccd1 _13159_/C sky130_fd_sc_hd__and2_1
XFILLER_124_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10266_ _18654_/Q _18076_/Q _19095_/Q _18999_/Q _09937_/S _10266_/S1 vssd1 vssd1
+ vccd1 vccd1 _10266_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1310 _11741_/A2 vssd1 vssd1 vccd1 vccd1 _11726_/B sky130_fd_sc_hd__buf_4
X_12005_ _17772_/Q _16540_/A0 _12022_/S vssd1 vssd1 vccd1 vccd1 _17772_/D sky130_fd_sc_hd__mux2_1
Xfanout1321 _09099_/Y vssd1 vssd1 vccd1 vccd1 _09106_/B sky130_fd_sc_hd__clkbuf_16
X_17862_ _17865_/CLK _17862_/D vssd1 vssd1 vccd1 vccd1 _17862_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1332 _10265_/A vssd1 vssd1 vccd1 vccd1 _10315_/S sky130_fd_sc_hd__buf_6
XFILLER_39_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1343 _10841_/C1 vssd1 vssd1 vccd1 vccd1 _10618_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10197_ _17917_/Q _11490_/B _11489_/B1 _10196_/Y vssd1 vssd1 vccd1 vccd1 _10233_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_238_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1354 _09919_/C1 vssd1 vssd1 vccd1 vccd1 _09914_/C1 sky130_fd_sc_hd__buf_4
X_19601_ _19601_/CLK _19601_/D vssd1 vssd1 vccd1 vccd1 _19601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16813_ _19293_/Q _16815_/C _16812_/Y vssd1 vssd1 vccd1 vccd1 _19293_/D sky130_fd_sc_hd__a21oi_1
XFILLER_213_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1365 _10856_/C vssd1 vssd1 vccd1 vccd1 _11325_/S sky130_fd_sc_hd__buf_6
Xfanout1376 _09843_/S vssd1 vssd1 vccd1 vccd1 _10634_/S0 sky130_fd_sc_hd__clkbuf_4
XFILLER_266_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17793_ _19650_/CLK _17793_/D vssd1 vssd1 vccd1 vccd1 _17793_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1387 _11147_/S vssd1 vssd1 vccd1 vccd1 _10001_/S sky130_fd_sc_hd__buf_6
XFILLER_282_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1398 fanout1407/X vssd1 vssd1 vccd1 vccd1 _10249_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_19_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19532_ _19533_/CLK _19532_/D vssd1 vssd1 vccd1 vccd1 _19532_/Q sky130_fd_sc_hd__dfxtp_1
X_16744_ _16752_/A _16744_/B _16746_/B vssd1 vssd1 vccd1 vccd1 _19267_/D sky130_fd_sc_hd__nor3_1
XFILLER_281_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13956_ _13758_/A _13941_/X _13956_/B1 vssd1 vssd1 vccd1 vccd1 _13956_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12907_ _17826_/Q _13942_/A2 _13942_/B1 _17858_/Q vssd1 vssd1 vccd1 vccd1 _12907_/X
+ sky130_fd_sc_hd__a22o_1
X_19463_ _19464_/CLK _19463_/D vssd1 vssd1 vccd1 vccd1 _19463_/Q sky130_fd_sc_hd__dfxtp_4
X_16675_ _16776_/A _16675_/B _16675_/C vssd1 vssd1 vccd1 vccd1 _19246_/D sky130_fd_sc_hd__nor3_1
X_13887_ _13929_/A1 _13886_/X _13874_/X vssd1 vssd1 vccd1 vccd1 _13887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_235_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18414_ _19591_/CLK _18414_/D vssd1 vssd1 vccd1 vccd1 _18414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15626_ _19447_/Q _15661_/B _17199_/A vssd1 vssd1 vccd1 vccd1 _15626_/X sky130_fd_sc_hd__o21a_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _12836_/Y _13316_/B _12838_/S vssd1 vssd1 vccd1 vccd1 _12838_/X sky130_fd_sc_hd__mux2_1
XFILLER_261_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19394_ _19526_/CLK _19394_/D vssd1 vssd1 vccd1 vccd1 _19394_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18345_ _19653_/A _18345_/D vssd1 vssd1 vccd1 vccd1 _18345_/Q sky130_fd_sc_hd__dfxtp_1
X_12769_ _19233_/Q _13495_/A2 _13495_/B1 _19265_/Q vssd1 vssd1 vccd1 vccd1 _12769_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ _15557_/A _15557_/B _15557_/C vssd1 vssd1 vccd1 vccd1 _15558_/B sky130_fd_sc_hd__or3_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_168_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19448_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14508_ _17710_/A0 _18358_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _18358_/D sky130_fd_sc_hd__mux2_1
XFILLER_202_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18276_ _18593_/CLK _18276_/D vssd1 vssd1 vccd1 vccd1 _18276_/Q sky130_fd_sc_hd__dfxtp_1
X_15488_ _18579_/Q _15512_/C vssd1 vssd1 vccd1 vccd1 _15488_/X sky130_fd_sc_hd__xor2_1
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17227_ _14714_/A _17157_/A _17404_/A _17256_/B vssd1 vssd1 vccd1 vccd1 _17227_/X
+ sky130_fd_sc_hd__o22a_1
Xinput20 core_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
Xinput31 core_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_2
X_14439_ _18578_/Q _17354_/A vssd1 vssd1 vccd1 vccd1 _18291_/D sky130_fd_sc_hd__and2_2
XFILLER_128_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 core_wb_error_i vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_2
Xinput53 dout0[19] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput64 dout0[29] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_2
X_17158_ _19404_/Q _17124_/B _17453_/A _17158_/B2 vssd1 vssd1 vccd1 vccd1 _17159_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xinput75 dout0[39] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput86 dout0[49] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput97 dout0[59] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16109_ _18757_/Q _16139_/B vssd1 vssd1 vccd1 vccd1 _16109_/Y sky130_fd_sc_hd__nand2_1
X_09980_ _11518_/B2 _09980_/A2 _09979_/X _09523_/A vssd1 vssd1 vccd1 vccd1 _09980_/Y
+ sky130_fd_sc_hd__a22oi_4
X_17089_ _19378_/Q _17115_/B vssd1 vssd1 vccd1 vccd1 _17089_/X sky130_fd_sc_hd__or2_1
XFILLER_115_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08931_ _08939_/A _08913_/X _11216_/A2 vssd1 vssd1 vccd1 vccd1 _08948_/A sky130_fd_sc_hd__a21oi_4
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ _18406_/Q _18405_/Q vssd1 vssd1 vccd1 vccd1 _11689_/A sky130_fd_sc_hd__nand2b_4
XFILLER_257_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09414_ _09412_/X _09413_/X _09429_/S vssd1 vssd1 vccd1 vccd1 _09414_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09345_ _11017_/A1 _19562_/Q _09344_/S _19594_/Q _10250_/S vssd1 vssd1 vccd1 vccd1
+ _09345_/X sky130_fd_sc_hd__o221a_1
XFILLER_200_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09276_ _11459_/B1 _09261_/X _09274_/X _09275_/X vssd1 vssd1 vccd1 vccd1 _09276_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_139_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10120_ _11452_/A _10119_/X _10089_/Y _11790_/B vssd1 vssd1 vccd1 vccd1 _10121_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_161_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10051_ _18048_/Q _10816_/A2 _10050_/X _11189_/A vssd1 vssd1 vccd1 vccd1 _10051_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _13810_/A _13861_/A vssd1 vssd1 vccd1 vccd1 _13810_/X sky130_fd_sc_hd__or2_1
XFILLER_263_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ _14992_/A1 _13251_/X _14973_/B1 _18636_/Q _14741_/B vssd1 vssd1 vccd1 vccd1
+ _14790_/X sky130_fd_sc_hd__a221o_1
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13741_ _11583_/A _13971_/A2 _13739_/Y _13740_/Y _13579_/A vssd1 vssd1 vccd1 vccd1
+ _13741_/X sky130_fd_sc_hd__a221o_4
X_10953_ _11352_/A1 _19637_/Q _18926_/Q _11340_/B2 vssd1 vssd1 vccd1 vccd1 _10953_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_272_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13672_ _13968_/A1 _13662_/X _13671_/X _13323_/B vssd1 vssd1 vccd1 vccd1 _13672_/X
+ sky130_fd_sc_hd__a22o_1
X_16460_ _17692_/A0 _19067_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _19067_/D sky130_fd_sc_hd__mux2_1
XFILLER_243_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10884_ _11594_/A1 _19119_/Q _19151_/Q _11613_/S vssd1 vssd1 vccd1 vccd1 _10884_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12623_ _12622_/A _13226_/A _13261_/A vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__a21o_1
X_15411_ _19438_/Q _15411_/B vssd1 vssd1 vccd1 vccd1 _15411_/X sky130_fd_sc_hd__or2_1
XFILLER_188_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16391_ _17690_/A0 _19002_/Q _16391_/S vssd1 vssd1 vccd1 vccd1 _19002_/D sky130_fd_sc_hd__mux2_1
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18130_ _19453_/CLK _18130_/D vssd1 vssd1 vccd1 vccd1 _18130_/Q sky130_fd_sc_hd__dfxtp_4
X_15342_ _18573_/Q _15342_/B vssd1 vssd1 vccd1 vccd1 _15342_/Y sky130_fd_sc_hd__nor2_1
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12554_ _12554_/A _12554_/B _12563_/B vssd1 vssd1 vccd1 vccd1 _12561_/B sky130_fd_sc_hd__or3_4
XFILLER_129_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ _11506_/A1 _18951_/Q _18216_/Q _10424_/S vssd1 vssd1 vccd1 vccd1 _11505_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18061_ _19079_/CLK _18061_/D vssd1 vssd1 vccd1 vccd1 _18061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15273_ _15731_/B1 _15272_/X _19432_/Q _15411_/B vssd1 vssd1 vccd1 vccd1 _15274_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_12485_ _12553_/A _12553_/B vssd1 vssd1 vccd1 vccd1 _12572_/A sky130_fd_sc_hd__nand2_1
XFILLER_200_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17012_ _17587_/A _17044_/A2 _17011_/X _17346_/A vssd1 vssd1 vccd1 vccd1 _19342_/D
+ sky130_fd_sc_hd__o211a_1
X_14224_ _14224_/A _14224_/B vssd1 vssd1 vccd1 vccd1 _14224_/Y sky130_fd_sc_hd__nand2_1
X_11436_ _11434_/X _11435_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _11436_/X sky130_fd_sc_hd__mux2_1
XFILLER_208_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14155_ _14155_/A _14155_/B vssd1 vssd1 vccd1 vccd1 _14155_/Y sky130_fd_sc_hd__nor2_1
X_11367_ _11368_/A _12596_/B vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__nor2_2
X_13106_ _19303_/Q _13952_/A2 _12551_/Y vssd1 vssd1 vccd1 vccd1 _13106_/X sky130_fd_sc_hd__a21o_1
X_10318_ _11173_/S _10316_/X _10317_/X vssd1 vssd1 vccd1 vccd1 _10318_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14086_ _17669_/A0 _18026_/Q _14106_/S vssd1 vssd1 vccd1 vccd1 _18026_/D sky130_fd_sc_hd__mux2_1
XFILLER_258_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18963_ _19155_/CLK _18963_/D vssd1 vssd1 vccd1 vccd1 _18963_/Q sky130_fd_sc_hd__dfxtp_1
X_11298_ _09987_/A _11297_/X _11295_/X vssd1 vssd1 vccd1 vccd1 _11298_/X sky130_fd_sc_hd__o21a_1
XFILLER_79_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17914_ _18881_/CLK _17914_/D vssd1 vssd1 vccd1 vccd1 _17914_/Q sky130_fd_sc_hd__dfxtp_4
X_13037_ _12803_/A _12826_/A _13089_/A vssd1 vssd1 vccd1 vccd1 _13038_/B sky130_fd_sc_hd__mux2_1
X_10249_ _18622_/Q _18193_/Q _10249_/S vssd1 vssd1 vccd1 vccd1 _10249_/X sky130_fd_sc_hd__mux2_1
X_18894_ _19632_/CLK _18894_/D vssd1 vssd1 vccd1 vccd1 _18894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1140 _09434_/X vssd1 vssd1 vccd1 vccd1 _09437_/B sky130_fd_sc_hd__buf_6
Xfanout1151 _09079_/Y vssd1 vssd1 vccd1 vccd1 _13421_/A sky130_fd_sc_hd__buf_6
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1162 _15954_/X vssd1 vssd1 vccd1 vccd1 _16003_/A2 sky130_fd_sc_hd__buf_4
X_17845_ _19470_/CLK _17845_/D vssd1 vssd1 vccd1 vccd1 _17845_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_78_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1173 _15946_/A2 vssd1 vssd1 vccd1 vccd1 _15943_/A2 sky130_fd_sc_hd__buf_4
XFILLER_226_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1184 _12317_/X vssd1 vssd1 vccd1 vccd1 _15526_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_282_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1195 _16893_/B1 vssd1 vssd1 vccd1 vccd1 _16969_/B1 sky130_fd_sc_hd__buf_4
XFILLER_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17776_ _19604_/CLK _17776_/D vssd1 vssd1 vccd1 vccd1 _17776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14988_ _14988_/A vssd1 vssd1 vccd1 vccd1 _14988_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_207_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19515_ _19546_/CLK _19515_/D vssd1 vssd1 vccd1 vccd1 _19515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16727_ _19261_/Q _16729_/C _19262_/Q vssd1 vssd1 vccd1 vccd1 _16730_/B sky130_fd_sc_hd__a21oi_1
X_13939_ _12442_/A _12448_/C _13937_/Y _13938_/Y _12762_/B vssd1 vssd1 vccd1 vccd1
+ _13939_/X sky130_fd_sc_hd__a221o_4
XFILLER_235_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19446_ _19546_/CLK _19446_/D vssd1 vssd1 vccd1 vccd1 _19446_/Q sky130_fd_sc_hd__dfxtp_1
X_16658_ _19241_/Q _19240_/Q _16658_/C vssd1 vssd1 vccd1 vccd1 _16664_/C sky130_fd_sc_hd__and3_1
XFILLER_250_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15609_ _19478_/Q _19412_/Q vssd1 vssd1 vccd1 vccd1 _15610_/B sky130_fd_sc_hd__nor2_1
X_19377_ _19506_/CLK _19377_/D vssd1 vssd1 vccd1 vccd1 _19377_/Q sky130_fd_sc_hd__dfxtp_2
X_16589_ _16622_/A0 _19193_/Q _16589_/S vssd1 vssd1 vccd1 vccd1 _19193_/D sky130_fd_sc_hd__mux2_1
XFILLER_222_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09130_ _18637_/Q _18059_/Q _09269_/S vssd1 vssd1 vccd1 vccd1 _09130_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18328_ _19575_/CLK _18328_/D vssd1 vssd1 vccd1 vccd1 _18328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_249_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09061_ _12665_/A _12264_/A vssd1 vssd1 vccd1 vccd1 _12756_/B sky130_fd_sc_hd__nor2_4
X_18259_ _19644_/CLK _18259_/D vssd1 vssd1 vccd1 vccd1 _18259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09963_ _09959_/X _09962_/X _10746_/S vssd1 vssd1 vccd1 vccd1 _09963_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_65_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19631_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08914_ _08932_/A _12051_/A _17802_/Q vssd1 vssd1 vccd1 vccd1 _08914_/X sky130_fd_sc_hd__or3b_4
XFILLER_98_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _11210_/A1 _16462_/A0 _09893_/Y _11055_/B2 vssd1 vssd1 vccd1 vccd1 _15130_/A
+ sky130_fd_sc_hd__o2bb2a_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08845_ _10027_/A vssd1 vssd1 vccd1 vccd1 _08845_/Y sky130_fd_sc_hd__inv_6
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_507 _17587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_518 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_529 _11853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09328_ _09039_/B _11141_/B _09327_/X vssd1 vssd1 vccd1 vccd1 _09328_/X sky130_fd_sc_hd__o21ba_1
XFILLER_179_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09259_ _09272_/A1 _19563_/Q _09269_/S _19595_/Q _09914_/C1 vssd1 vssd1 vccd1 vccd1
+ _09259_/X sky130_fd_sc_hd__o221a_1
XFILLER_167_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12270_ _12271_/A _12271_/B vssd1 vssd1 vccd1 vccd1 _15835_/B sky130_fd_sc_hd__nor2_2
XFILLER_119_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11221_ _09050_/X _11217_/X _11219_/Y _11220_/X vssd1 vssd1 vccd1 vccd1 _11221_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_175_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11152_ _18548_/Q _11226_/S vssd1 vssd1 vccd1 vccd1 _11152_/X sky130_fd_sc_hd__or2_1
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10103_ _10253_/A _18809_/Q _10176_/S vssd1 vssd1 vccd1 vccd1 _10103_/X sky130_fd_sc_hd__and3_1
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15960_ _18695_/Q _15970_/A2 _15976_/B1 _18744_/Q _15976_/C1 vssd1 vssd1 vccd1 vccd1
+ _15960_/X sky130_fd_sc_hd__a221o_1
X_11083_ _19635_/Q _18924_/Q _11094_/S vssd1 vssd1 vccd1 vccd1 _11083_/X sky130_fd_sc_hd__mux2_1
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput210 localMemory_wb_adr_i[6] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput221 localMemory_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input221/X sky130_fd_sc_hd__clkbuf_16
XFILLER_68_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput232 localMemory_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 input232/X sky130_fd_sc_hd__buf_12
X_14911_ _17812_/Q _14911_/B vssd1 vssd1 vccd1 vccd1 _14911_/X sky130_fd_sc_hd__or2_1
X_10034_ _18843_/Q _18875_/Q _10496_/B vssd1 vssd1 vccd1 vccd1 _10034_/X sky130_fd_sc_hd__mux2_1
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput243 localMemory_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input243/X sky130_fd_sc_hd__buf_8
XFILLER_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput254 manufacturerID[10] vssd1 vssd1 vccd1 vccd1 _15887_/A sky130_fd_sc_hd__buf_4
X_15891_ _18672_/Q _15906_/A2 _15903_/B1 _15890_/X vssd1 vssd1 vccd1 vccd1 _15891_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput265 partID[10] vssd1 vssd1 vccd1 vccd1 _15920_/A sky130_fd_sc_hd__buf_2
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput276 partID[6] vssd1 vssd1 vccd1 vccd1 _15908_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_263_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17630_ _17663_/A0 _19558_/Q _17654_/S vssd1 vssd1 vccd1 vccd1 _19558_/D sky130_fd_sc_hd__mux2_1
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _18116_/Q _14994_/B _14771_/X _14841_/X vssd1 vssd1 vccd1 vccd1 _14842_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17561_ _19523_/Q _17561_/B vssd1 vssd1 vccd1 vccd1 _17561_/X sky130_fd_sc_hd__or2_1
X_11985_ _12460_/A _14487_/A _11985_/C _09055_/B vssd1 vssd1 vccd1 vccd1 _16459_/B
+ sky130_fd_sc_hd__or4b_4
X_14773_ _14865_/A1 _14772_/X _14865_/B1 vssd1 vssd1 vccd1 vccd1 _14773_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19300_ _19300_/CLK _19300_/D vssd1 vssd1 vccd1 vccd1 _19300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16512_ _16545_/A0 _19118_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _19118_/D sky130_fd_sc_hd__mux2_1
X_13724_ _13929_/A1 _13723_/X _13711_/Y vssd1 vssd1 vccd1 vccd1 _13724_/Y sky130_fd_sc_hd__a21oi_1
X_10936_ _18830_/Q _11300_/B vssd1 vssd1 vccd1 vccd1 _10936_/X sky130_fd_sc_hd__or2_1
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17492_ _18121_/Q _17539_/C1 _17490_/X _17491_/X vssd1 vssd1 vccd1 vccd1 _17492_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19231_ _19231_/CLK _19231_/D vssd1 vssd1 vccd1 vccd1 _19231_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_140_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16443_ _19051_/Q _16542_/A0 _16454_/S vssd1 vssd1 vccd1 vccd1 _19051_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10867_ _10861_/X _10863_/X _10866_/X _11578_/S _11588_/B1 vssd1 vssd1 vccd1 vccd1
+ _10867_/X sky130_fd_sc_hd__o221a_1
X_13655_ _19446_/Q _13655_/A2 _13653_/X _13654_/X _13655_/C1 vssd1 vssd1 vccd1 vccd1
+ _13655_/X sky130_fd_sc_hd__o221a_1
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _12900_/A _12900_/B _12602_/X vssd1 vssd1 vccd1 vccd1 _12957_/B sky130_fd_sc_hd__o21a_2
X_19162_ _19163_/CLK _19162_/D vssd1 vssd1 vccd1 vccd1 _19162_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _19542_/Q _13946_/B vssd1 vssd1 vccd1 vccd1 _13586_/X sky130_fd_sc_hd__or2_1
X_16374_ _16507_/A0 _18985_/Q _16391_/S vssd1 vssd1 vccd1 vccd1 _18985_/D sky130_fd_sc_hd__mux2_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _11596_/A1 _19575_/Q _11604_/S _19607_/Q _11355_/A1 vssd1 vssd1 vccd1 vccd1
+ _10798_/X sky130_fd_sc_hd__o221a_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _19448_/CLK _18113_/D vssd1 vssd1 vccd1 vccd1 _18113_/Q sky130_fd_sc_hd__dfxtp_4
X_12537_ _12576_/A _12552_/B vssd1 vssd1 vccd1 vccd1 _12538_/B sky130_fd_sc_hd__or2_4
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15325_ _19466_/Q _15324_/X _15400_/S vssd1 vssd1 vccd1 vccd1 _15325_/X sky130_fd_sc_hd__mux2_1
X_19093_ _19157_/CLK _19093_/D vssd1 vssd1 vccd1 vccd1 _19093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ _19614_/CLK _18044_/D vssd1 vssd1 vccd1 vccd1 _18044_/Q sky130_fd_sc_hd__dfxtp_1
X_12468_ _16852_/A _12468_/B vssd1 vssd1 vccd1 vccd1 _12468_/Y sky130_fd_sc_hd__nand2_2
X_15256_ _17389_/B1 _15255_/X _15424_/C1 vssd1 vssd1 vccd1 vccd1 _15256_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11419_ _18856_/Q _18888_/Q _19048_/Q _19016_/Q _09290_/S _11503_/S1 vssd1 vssd1
+ vccd1 vccd1 _11419_/X sky130_fd_sc_hd__mux4_1
X_14207_ _18275_/Q _14247_/A2 _14206_/X _17380_/A vssd1 vssd1 vccd1 vccd1 _18101_/D
+ sky130_fd_sc_hd__o211a_1
X_15187_ _19460_/Q _19394_/Q vssd1 vssd1 vccd1 vccd1 _15188_/B sky130_fd_sc_hd__nand2_1
X_12399_ _12429_/A1 _09236_/A _09657_/X _12417_/B1 _18393_/Q vssd1 vssd1 vccd1 vccd1
+ _12400_/B sky130_fd_sc_hd__o32ai_2
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ _16522_/A0 _18077_/Q _14139_/S vssd1 vssd1 vccd1 vccd1 _18077_/D sky130_fd_sc_hd__mux2_1
XFILLER_235_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14069_ _16553_/A0 _18011_/Q _14072_/S vssd1 vssd1 vccd1 vccd1 _18011_/D sky130_fd_sc_hd__mux2_1
X_18946_ _19614_/CLK _18946_/D vssd1 vssd1 vccd1 vccd1 _18946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18877_ _19133_/CLK _18877_/D vssd1 vssd1 vccd1 vccd1 _18877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17828_ _18761_/CLK _17828_/D vssd1 vssd1 vccd1 vccd1 _17828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17759_ _19047_/CLK _17759_/D vssd1 vssd1 vccd1 vccd1 _17759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_183_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17931_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_112_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19280_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_222_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19429_ _19526_/CLK _19429_/D vssd1 vssd1 vccd1 vccd1 _19429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09113_ _18543_/Q _11455_/S vssd1 vssd1 vccd1 vccd1 _09113_/X sky130_fd_sc_hd__or2_1
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09044_ input109/X input144/X _09651_/S vssd1 vssd1 vccd1 vccd1 _09045_/B sky130_fd_sc_hd__mux2_4
XFILLER_276_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout900 _16204_/A0 vssd1 vssd1 vccd1 vccd1 _17701_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout1909 _11712_/A vssd1 vssd1 vccd1 vccd1 _14846_/B1 sky130_fd_sc_hd__buf_4
Xfanout911 _16393_/Y vssd1 vssd1 vccd1 vccd1 _16425_/S sky130_fd_sc_hd__buf_12
XFILLER_104_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout922 _16245_/S vssd1 vssd1 vccd1 vccd1 _16255_/S sky130_fd_sc_hd__buf_12
X_09946_ _09944_/X _09945_/Y _09946_/B1 vssd1 vssd1 vccd1 vccd1 _09946_/X sky130_fd_sc_hd__a21o_1
Xfanout933 _14983_/B1 vssd1 vssd1 vccd1 vccd1 _15003_/B1 sky130_fd_sc_hd__buf_4
Xfanout944 _14671_/X vssd1 vssd1 vccd1 vccd1 _14994_/B sky130_fd_sc_hd__buf_4
Xfanout955 _14628_/S vssd1 vssd1 vccd1 vccd1 _14630_/S sky130_fd_sc_hd__buf_12
XFILLER_258_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout966 _14075_/Y vssd1 vssd1 vccd1 vccd1 _14098_/S sky130_fd_sc_hd__buf_6
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout977 _12463_/X vssd1 vssd1 vccd1 vccd1 _13527_/B1 sky130_fd_sc_hd__buf_4
XFILLER_218_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _09877_/A _09877_/B vssd1 vssd1 vccd1 vccd1 _09877_/Y sky130_fd_sc_hd__nor2_1
XFILLER_245_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout988 _12449_/X vssd1 vssd1 vccd1 vccd1 _13973_/A2 sky130_fd_sc_hd__buf_6
XFILLER_86_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout999 _10459_/X vssd1 vssd1 vccd1 vccd1 _17684_/A0 sky130_fd_sc_hd__buf_4
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _08828_/A vssd1 vssd1 vccd1 vccd1 _08828_/Y sky130_fd_sc_hd__inv_2
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_304 _18113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_315 _18102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 _11953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_337 _10194_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_348 _10211_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11770_ _18588_/Q _14349_/B _11770_/B1 _13807_/B vssd1 vssd1 vccd1 vccd1 _11770_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_359 _15549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10721_ _18038_/Q _18006_/Q _10721_/S vssd1 vssd1 vccd1 vccd1 _10721_/X sky130_fd_sc_hd__mux2_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13968_/A1 _13421_/Y _13439_/X _13420_/X _13968_/B2 vssd1 vssd1 vccd1 vccd1
+ _13440_/X sky130_fd_sc_hd__a32o_1
X_10652_ _10643_/S _10650_/X _10651_/X _10653_/C1 vssd1 vssd1 vccd1 vccd1 _10652_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13371_ _19246_/Q _13425_/A2 _13425_/B1 _19278_/Q vssd1 vssd1 vccd1 vccd1 _13371_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10583_ _19059_/Q _19027_/Q _10656_/S vssd1 vssd1 vccd1 vccd1 _10583_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15110_ _15111_/A _15133_/B vssd1 vssd1 vccd1 vccd1 _15110_/X sky130_fd_sc_hd__and2_2
X_12322_ _12323_/A _12323_/B vssd1 vssd1 vccd1 vccd1 _12322_/Y sky130_fd_sc_hd__nor2_8
X_16090_ _16096_/A1 _16089_/Y _17725_/C1 vssd1 vssd1 vccd1 vccd1 _18747_/D sky130_fd_sc_hd__a21oi_1
XFILLER_194_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15041_ _15013_/A _15013_/B input252/X _11711_/A vssd1 vssd1 vccd1 vccd1 _15043_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12253_ _17883_/Q _17884_/Q _12253_/C vssd1 vssd1 vccd1 vccd1 _12256_/B sky130_fd_sc_hd__and3_1
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ _11618_/A1 _18323_/Q _17774_/Q _10726_/S vssd1 vssd1 vccd1 vccd1 _11204_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12184_ _17857_/Q _17858_/Q _12184_/C vssd1 vssd1 vccd1 vccd1 _12186_/B sky130_fd_sc_hd__and3_1
XFILLER_122_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18800_ _19607_/CLK _18800_/D vssd1 vssd1 vccd1 vccd1 _18800_/Q sky130_fd_sc_hd__dfxtp_1
X_11135_ _18118_/Q _11134_/Y _11135_/S vssd1 vssd1 vccd1 vccd1 _11138_/B sky130_fd_sc_hd__mux2_2
XFILLER_96_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16992_ _17567_/A _17008_/A2 _16991_/X _17419_/C1 vssd1 vssd1 vccd1 vccd1 _19332_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ _18734_/CLK _18731_/D vssd1 vssd1 vccd1 vccd1 _18731_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_283_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15943_ _18690_/Q _15943_/A2 _15942_/X _15946_/C1 vssd1 vssd1 vccd1 vccd1 _18690_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11066_ _11066_/A _11066_/B vssd1 vssd1 vccd1 vccd1 _11066_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ _18843_/Q _18875_/Q _19035_/Q _19003_/Q _11070_/S _12320_/A vssd1 vssd1 vccd1
+ vccd1 _10017_/X sky130_fd_sc_hd__mux4_1
X_18662_ _18715_/CLK _18662_/D vssd1 vssd1 vccd1 vccd1 _18662_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _18667_/Q _15949_/A2 _15872_/X _15873_/X _15904_/C1 vssd1 vssd1 vccd1 vccd1
+ _18667_/D sky130_fd_sc_hd__o221a_1
XFILLER_264_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17613_ _19488_/Q _15093_/D _17556_/A _17199_/B _17556_/X vssd1 vssd1 vccd1 vccd1
+ _17613_/X sky130_fd_sc_hd__a221o_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _14825_/A vssd1 vssd1 vccd1 vccd1 _14825_/Y sky130_fd_sc_hd__inv_2
XFILLER_218_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _18593_/CLK _18593_/D vssd1 vssd1 vccd1 vccd1 _18593_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17544_ _17544_/A _17544_/B vssd1 vssd1 vccd1 vccd1 _17544_/X sky130_fd_sc_hd__and2_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _14718_/A _14755_/X _14846_/B1 vssd1 vssd1 vccd1 vccd1 _14756_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_204_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11968_ _18514_/Q _11720_/X _11918_/X _11968_/B2 vssd1 vssd1 vccd1 vccd1 _11968_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13707_ _15133_/A _13703_/X _13706_/X _13869_/B2 vssd1 vssd1 vccd1 vccd1 _13707_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10919_ _11305_/A1 _19150_/Q _11094_/S _19118_/Q _11562_/S vssd1 vssd1 vccd1 vccd1
+ _10919_/X sky130_fd_sc_hd__o221a_1
X_17475_ _13512_/B _17475_/A2 _17475_/B1 _17807_/Q _17550_/A vssd1 vssd1 vccd1 vccd1
+ _17475_/X sky130_fd_sc_hd__a221o_1
XFILLER_205_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14687_ _14687_/A _14687_/B vssd1 vssd1 vccd1 vccd1 _14688_/D sky130_fd_sc_hd__or2_1
X_11899_ _11899_/A _11899_/B _11899_/C vssd1 vssd1 vccd1 vccd1 _11899_/X sky130_fd_sc_hd__and3_4
XFILLER_260_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19214_ _19637_/CLK _19214_/D vssd1 vssd1 vccd1 vccd1 _19214_/Q sky130_fd_sc_hd__dfxtp_1
X_16426_ _16426_/A _16591_/B vssd1 vssd1 vccd1 vccd1 _16426_/X sky130_fd_sc_hd__and2_1
X_13638_ _13758_/A _13638_/B vssd1 vssd1 vccd1 vccd1 _13638_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19145_ _19600_/CLK _19145_/D vssd1 vssd1 vccd1 vccd1 _19145_/Q sky130_fd_sc_hd__dfxtp_1
X_16357_ _18969_/Q _16490_/A0 _16357_/S vssd1 vssd1 vccd1 vccd1 _18969_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13569_ _13861_/A _14148_/A _13892_/B1 vssd1 vssd1 vccd1 vccd1 _13569_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15308_ _15306_/Y _15308_/B vssd1 vssd1 vccd1 vccd1 _15365_/C sky130_fd_sc_hd__and2b_1
X_19076_ _19076_/CLK _19076_/D vssd1 vssd1 vccd1 vccd1 _19076_/Q sky130_fd_sc_hd__dfxtp_1
X_16288_ _17719_/A0 _18902_/Q _16288_/S vssd1 vssd1 vccd1 vccd1 _18902_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18027_ _18543_/CLK _18027_/D vssd1 vssd1 vccd1 vccd1 _18027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15239_ _15304_/A1 _13122_/Y _15285_/A3 _15238_/X vssd1 vssd1 vccd1 vccd1 _15239_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_259_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09800_ _11284_/A1 _19557_/Q _09797_/S _19589_/Q _10040_/S vssd1 vssd1 vccd1 vccd1
+ _09800_/X sky130_fd_sc_hd__o221a_1
XFILLER_259_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09731_ _11518_/B2 _09662_/X _09730_/X _09523_/A vssd1 vssd1 vccd1 vccd1 _15173_/A
+ sky130_fd_sc_hd__a22o_4
X_18929_ _19640_/CLK _18929_/D vssd1 vssd1 vccd1 vccd1 _18929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_268_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09662_ _17956_/Q _11216_/A2 _08947_/X _17924_/Q _09661_/X vssd1 vssd1 vccd1 vccd1
+ _09662_/X sky130_fd_sc_hd__a221o_4
XFILLER_55_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09593_ _18312_/Q _17763_/Q _10362_/S vssd1 vssd1 vccd1 vccd1 _09593_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19587_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09027_ _09027_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _11219_/A sky130_fd_sc_hd__nand2_2
XFILLER_237_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1706 _09350_/S vssd1 vssd1 vccd1 vccd1 _09264_/S sky130_fd_sc_hd__buf_12
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1717 _16898_/A1 vssd1 vssd1 vccd1 vccd1 _16970_/A1 sky130_fd_sc_hd__buf_8
Xfanout730 _11451_/X vssd1 vssd1 vccd1 vccd1 _16538_/A0 sky130_fd_sc_hd__buf_2
Xfanout1728 _08828_/A vssd1 vssd1 vccd1 vccd1 _16969_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout741 _17641_/A0 vssd1 vssd1 vccd1 vccd1 _16607_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_132_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1739 _15009_/A1 vssd1 vssd1 vccd1 vccd1 _14979_/A1 sky130_fd_sc_hd__buf_4
XFILLER_59_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09929_ _18844_/Q _11167_/B _09928_/X vssd1 vssd1 vccd1 vccd1 _09929_/X sky130_fd_sc_hd__a21o_1
Xfanout752 _13390_/S vssd1 vssd1 vccd1 vccd1 _13194_/S sky130_fd_sc_hd__buf_4
Xfanout763 _09054_/X vssd1 vssd1 vccd1 vccd1 _16471_/A0 sky130_fd_sc_hd__buf_2
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout774 _17625_/Y vssd1 vssd1 vccd1 vccd1 _17648_/S sky130_fd_sc_hd__buf_6
XFILLER_246_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout785 _16525_/Y vssd1 vssd1 vccd1 vccd1 _16557_/S sky130_fd_sc_hd__buf_12
Xfanout796 _16326_/Y vssd1 vssd1 vccd1 vccd1 _16355_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_246_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12940_ _12800_/X _12824_/Y _12942_/S vssd1 vssd1 vccd1 vccd1 _13130_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _13079_/A _12866_/Y _12867_/X _12870_/X vssd1 vssd1 vccd1 vccd1 _12871_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_218_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _15450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _11780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ _17669_/A0 _18417_/Q _14630_/S vssd1 vssd1 vccd1 vccd1 _18417_/D sky130_fd_sc_hd__mux2_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_123 _11825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _11814_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11822_ _11844_/A _11822_/B vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__and2_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15590_/A _15590_/B vssd1 vssd1 vccd1 vccd1 _15591_/B sky130_fd_sc_hd__nor2_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _11868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _11872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _13049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_178 _13444_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11753_ _13225_/A _11753_/B vssd1 vssd1 vccd1 vccd1 _13224_/A sky130_fd_sc_hd__xor2_4
X_14541_ _18379_/Q _14559_/A2 _14559_/B1 input38/X vssd1 vssd1 vccd1 vccd1 _14542_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _13723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _11250_/A1 _18226_/Q _11154_/S _18961_/Q vssd1 vssd1 vccd1 vccd1 _10704_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_241_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17260_ _19437_/Q _17310_/B _17259_/X vssd1 vssd1 vccd1 vccd1 _17261_/B sky130_fd_sc_hd__a21oi_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ _18324_/Q _17676_/A0 _14486_/S vssd1 vssd1 vccd1 vccd1 _18324_/D sky130_fd_sc_hd__mux2_1
X_11684_ _13476_/B _13443_/B _13402_/B _11684_/D vssd1 vssd1 vccd1 vccd1 _11685_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_201_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16211_ _16608_/A0 _18827_/Q _16222_/S vssd1 vssd1 vccd1 vccd1 _18827_/D sky130_fd_sc_hd__mux2_1
X_13423_ _17838_/Q _13844_/A2 _13844_/B1 _17870_/Q vssd1 vssd1 vccd1 vccd1 _13423_/X
+ sky130_fd_sc_hd__a22o_1
X_10635_ _10618_/S _10634_/X _09106_/B vssd1 vssd1 vccd1 vccd1 _10635_/X sky130_fd_sc_hd__o21a_1
XFILLER_139_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17191_ _19415_/Q fanout533/X _17508_/A _17119_/B vssd1 vssd1 vccd1 vccd1 _17192_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16142_ _16142_/A1 _16141_/Y _16142_/B1 vssd1 vssd1 vccd1 vccd1 _18773_/D sky130_fd_sc_hd__a21oi_1
XFILLER_220_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13354_ _13354_/A _13354_/B vssd1 vssd1 vccd1 vccd1 _13354_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10566_ _18331_/Q _17782_/Q _10645_/S vssd1 vssd1 vccd1 vccd1 _10566_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12305_ _18097_/Q _12305_/A2 _12305_/B1 _18520_/Q vssd1 vssd1 vccd1 vccd1 _14687_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13285_ _17834_/Q _13944_/B _13284_/X vssd1 vssd1 vccd1 vccd1 _13285_/X sky130_fd_sc_hd__o21a_1
XFILLER_182_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16073_ _16020_/A _18740_/Q _14427_/B _16072_/Y vssd1 vssd1 vccd1 vccd1 _18740_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10497_ _18073_/Q _10816_/A2 _10496_/X _11189_/A vssd1 vssd1 vccd1 vccd1 _10497_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15024_ _18513_/Q input213/X _15024_/S vssd1 vssd1 vccd1 vccd1 _18513_/D sky130_fd_sc_hd__mux2_1
X_12236_ _17877_/Q _12234_/B _12235_/Y vssd1 vssd1 vccd1 vccd1 _17877_/D sky130_fd_sc_hd__o21a_1
XFILLER_154_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12167_ _17851_/Q _12168_/C _17852_/Q vssd1 vssd1 vccd1 vccd1 _12169_/B sky130_fd_sc_hd__a21oi_1
XFILLER_2_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11118_ _11352_/A1 _19212_/Q _19180_/Q _11125_/B2 vssd1 vssd1 vccd1 vccd1 _11118_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12098_ _12107_/A _12098_/B vssd1 vssd1 vccd1 vccd1 _12098_/Y sky130_fd_sc_hd__nor2_1
X_16975_ _17052_/A _16975_/B _16975_/C vssd1 vssd1 vccd1 vccd1 _17047_/B sky130_fd_sc_hd__or3_2
XFILLER_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18714_ _18715_/CLK _18714_/D vssd1 vssd1 vccd1 vccd1 _18714_/Q sky130_fd_sc_hd__dfxtp_1
X_15926_ input1/X input267/X _15947_/S vssd1 vssd1 vccd1 vccd1 _15926_/X sky130_fd_sc_hd__mux2_1
X_11049_ _11047_/X _11048_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _11049_/X sky130_fd_sc_hd__mux2_1
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 coreIndex[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_6
XFILLER_265_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18645_ _19114_/CLK _18645_/D vssd1 vssd1 vccd1 vccd1 _18645_/Q sky130_fd_sc_hd__dfxtp_4
X_15857_ _15857_/A _15881_/B _15908_/C vssd1 vssd1 vccd1 vccd1 _15857_/X sky130_fd_sc_hd__and3_1
XFILLER_252_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14808_ _18482_/Q _15001_/A2 _14807_/Y _12249_/A vssd1 vssd1 vccd1 vccd1 _18482_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18576_ _19537_/CLK _18576_/D vssd1 vssd1 vccd1 vccd1 _18576_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _15788_/A _15788_/B vssd1 vssd1 vccd1 vccd1 _15788_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_212_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17527_ _17527_/A1 _17525_/X _17526_/Y _17545_/C1 vssd1 vssd1 vccd1 vccd1 _17527_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_205_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14739_ _14736_/Y _14738_/Y _14879_/B1 vssd1 vssd1 vccd1 vccd1 _14739_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17458_ _18114_/Q _17463_/A2 _17456_/X _17457_/Y vssd1 vssd1 vccd1 vccd1 _17458_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16409_ _16607_/A0 _19018_/Q _16420_/S vssd1 vssd1 vccd1 vccd1 _19018_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17389_ _17118_/B _16973_/B _16979_/Y _17389_/B1 vssd1 vssd1 vccd1 vccd1 _17389_/X
+ sky130_fd_sc_hd__a31o_1
X_19128_ _19613_/CLK _19128_/D vssd1 vssd1 vccd1 vccd1 _19128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19059_ _19638_/CLK _19059_/D vssd1 vssd1 vccd1 vccd1 _19059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput300 _11916_/X vssd1 vssd1 vccd1 vccd1 addr1[6] sky130_fd_sc_hd__buf_4
XFILLER_134_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput311 _11759_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[15] sky130_fd_sc_hd__buf_4
XFILLER_145_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput322 _11769_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[25] sky130_fd_sc_hd__buf_4
Xoutput333 _08884_/X vssd1 vssd1 vccd1 vccd1 core_wb_cyc_o sky130_fd_sc_hd__buf_4
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput344 _11853_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[19] sky130_fd_sc_hd__buf_4
XFILLER_160_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput355 _11899_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[29] sky130_fd_sc_hd__buf_4
XFILLER_273_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput366 _11772_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[0] sky130_fd_sc_hd__buf_4
Xoutput377 _11930_/X vssd1 vssd1 vccd1 vccd1 din0[10] sky130_fd_sc_hd__buf_4
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput388 _11940_/X vssd1 vssd1 vccd1 vccd1 din0[20] sky130_fd_sc_hd__buf_4
Xoutput399 _11950_/X vssd1 vssd1 vccd1 vccd1 din0[30] sky130_fd_sc_hd__buf_4
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09714_ _09710_/X _09713_/X _10746_/S vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__mux2_1
XFILLER_262_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ _12614_/B _09647_/B vssd1 vssd1 vccd1 vccd1 _13044_/S sky130_fd_sc_hd__and2_2
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09576_ _17957_/Q _11216_/A2 _08947_/X _17925_/Q _09575_/X vssd1 vssd1 vccd1 vccd1
+ _09611_/B sky130_fd_sc_hd__a221o_4
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_169_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ _11513_/A1 _19580_/Q _10424_/S _19612_/Q _10427_/C1 vssd1 vssd1 vccd1 vccd1
+ _10420_/X sky130_fd_sc_hd__o221a_1
XFILLER_137_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10351_ _19126_/Q _19158_/Q _10353_/S vssd1 vssd1 vccd1 vccd1 _10351_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13070_ _19302_/Q _13174_/A _13068_/X _13069_/X _12551_/Y vssd1 vssd1 vccd1 vccd1
+ _13070_/X sky130_fd_sc_hd__a221o_2
XFILLER_279_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10282_ _10282_/A1 _18232_/Q _10281_/S _18967_/Q _10300_/S vssd1 vssd1 vccd1 vccd1
+ _10282_/X sky130_fd_sc_hd__o221a_1
XFILLER_183_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12021_ _17788_/Q _17722_/A0 _12021_/S vssd1 vssd1 vccd1 vccd1 _17788_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1503 _08968_/S0 vssd1 vssd1 vccd1 vccd1 _09952_/S sky130_fd_sc_hd__buf_6
XFILLER_160_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1514 fanout1524/X vssd1 vssd1 vccd1 vccd1 fanout1514/X sky130_fd_sc_hd__clkbuf_8
Xfanout1525 _08901_/Y vssd1 vssd1 vccd1 vccd1 fanout1525/X sky130_fd_sc_hd__buf_12
Xfanout1536 _10346_/S vssd1 vssd1 vccd1 vccd1 _10200_/S sky130_fd_sc_hd__buf_6
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1547 _11616_/S vssd1 vssd1 vccd1 vccd1 _10745_/S sky130_fd_sc_hd__buf_6
XFILLER_265_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout560 _15537_/B1 vssd1 vssd1 vccd1 vccd1 _15690_/A sky130_fd_sc_hd__buf_2
XFILLER_59_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1558 _09374_/S vssd1 vssd1 vccd1 vccd1 _10427_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout1569 _11508_/B1 vssd1 vssd1 vccd1 vccd1 _11495_/B1 sky130_fd_sc_hd__buf_12
Xfanout571 _15381_/A3 vssd1 vssd1 vccd1 vccd1 _15285_/A3 sky130_fd_sc_hd__buf_6
X_16760_ _16768_/A _16760_/B _16762_/B vssd1 vssd1 vccd1 vccd1 _19273_/D sky130_fd_sc_hd__nor3_1
Xfanout582 _12338_/Y vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout593 _14247_/A2 vssd1 vssd1 vccd1 vccd1 _14261_/A2 sky130_fd_sc_hd__buf_4
XFILLER_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13972_ _13545_/A _13958_/A _13970_/X vssd1 vssd1 vccd1 vccd1 _13972_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_265_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15711_ _19483_/Q _19417_/Q vssd1 vssd1 vccd1 vccd1 _15713_/A sky130_fd_sc_hd__or2_1
XFILLER_262_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12923_ _13757_/A _13980_/B _12906_/X vssd1 vssd1 vccd1 vccd1 _12923_/Y sky130_fd_sc_hd__o21ai_1
X_16691_ _19249_/Q _16686_/B _16689_/Y vssd1 vssd1 vccd1 vccd1 _19249_/D sky130_fd_sc_hd__o21a_1
XFILLER_46_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18430_ _19154_/CLK _18430_/D vssd1 vssd1 vccd1 vccd1 _18430_/Q sky130_fd_sc_hd__dfxtp_1
X_15642_ _15558_/A _15558_/B _15638_/X _15641_/X vssd1 vssd1 vccd1 vccd1 _15644_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_73_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12854_ _19426_/Q _12582_/X _12578_/Y vssd1 vssd1 vccd1 vccd1 _12854_/X sky130_fd_sc_hd__o21ba_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _19216_/CLK _18361_/D vssd1 vssd1 vccd1 vccd1 _18361_/Q sky130_fd_sc_hd__dfxtp_1
X_11805_ _11820_/A _11804_/X _11803_/Y vssd1 vssd1 vccd1 vccd1 _11806_/C sky130_fd_sc_hd__a21oi_4
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15573_ _18582_/Q _15800_/A2 _15565_/Y _15572_/X _17376_/A vssd1 vssd1 vccd1 vccd1
+ _18582_/D sky130_fd_sc_hd__o221a_1
XFILLER_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _13438_/A _12766_/X _13956_/B1 vssd1 vssd1 vccd1 vccd1 _12785_/X sky130_fd_sc_hd__a21o_1
XFILLER_214_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _17310_/Y _17311_/X _17231_/A vssd1 vssd1 vccd1 vccd1 _19454_/D sky130_fd_sc_hd__a21oi_1
X_14524_ input42/X _08884_/X _17198_/A vssd1 vssd1 vccd1 vccd1 _14524_/X sky130_fd_sc_hd__a21o_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18292_ _18593_/CLK _18292_/D vssd1 vssd1 vccd1 vccd1 _18292_/Q sky130_fd_sc_hd__dfxtp_1
X_11736_ _18565_/Q _11741_/A2 _11769_/B1 _12956_/A vssd1 vssd1 vccd1 vccd1 _11736_/X
+ sky130_fd_sc_hd__a22o_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17243_ _17241_/Y _17242_/X _17255_/A vssd1 vssd1 vccd1 vccd1 _19431_/D sky130_fd_sc_hd__a21oi_1
XFILLER_186_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14455_ _18307_/Q _16526_/A0 _14477_/S vssd1 vssd1 vccd1 vccd1 _18307_/D sky130_fd_sc_hd__mux2_1
XFILLER_175_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ _11667_/A _13697_/A vssd1 vssd1 vccd1 vccd1 _13695_/A sky130_fd_sc_hd__xnor2_4
XFILLER_128_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13406_ _18116_/Q _13406_/B vssd1 vssd1 vccd1 vccd1 _13407_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10618_ _10616_/X _10617_/X _10618_/S vssd1 vssd1 vccd1 vccd1 _10618_/X sky130_fd_sc_hd__mux2_1
X_17174_ _17231_/A _17174_/B vssd1 vssd1 vccd1 vccd1 _19409_/D sky130_fd_sc_hd__nor2_1
X_14386_ _17693_/A0 _18237_/Q _14412_/S vssd1 vssd1 vccd1 vccd1 _18237_/D sky130_fd_sc_hd__mux2_1
X_11598_ _18625_/Q _18196_/Q _11598_/S vssd1 vssd1 vccd1 vccd1 _11598_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16125_ _18765_/Q _16139_/B vssd1 vssd1 vccd1 vccd1 _16125_/Y sky130_fd_sc_hd__nand2_1
X_10549_ _18556_/Q _18431_/Q _18040_/Q _18008_/Q _09108_/B _11559_/S1 vssd1 vssd1
+ vccd1 vccd1 _10549_/X sky130_fd_sc_hd__mux4_1
X_13337_ _19405_/Q _12579_/Y _12771_/X _13336_/X _12581_/Y vssd1 vssd1 vccd1 vccd1
+ _13337_/X sky130_fd_sc_hd__a221o_1
XFILLER_128_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16056_ _16075_/A _16056_/B vssd1 vssd1 vccd1 vccd1 _16056_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13268_ _13267_/A _13797_/A0 _13267_/Y _13358_/A1 vssd1 vssd1 vccd1 vccd1 _13268_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15007_ input67/X input102/X _15007_/S vssd1 vssd1 vccd1 vccd1 _15008_/A sky130_fd_sc_hd__mux2_2
X_12219_ _12219_/A _12224_/C vssd1 vssd1 vccd1 vccd1 _12219_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13199_ _13191_/X _13198_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _13199_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16958_ _16970_/A1 _17948_/Q _16957_/X vssd1 vssd1 vccd1 vccd1 _17205_/B sky130_fd_sc_hd__o21a_4
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15909_ _18678_/Q _15918_/A2 _15945_/C1 _15908_/X vssd1 vssd1 vccd1 vccd1 _15909_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16889_ _18753_/Q _16893_/A2 _16893_/B1 input217/X _12483_/A vssd1 vssd1 vccd1 vccd1
+ _16889_/X sky130_fd_sc_hd__a221o_1
XFILLER_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09430_ _10300_/S _09429_/X _08903_/A vssd1 vssd1 vccd1 vccd1 _09430_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18628_ _18632_/CLK _18628_/D vssd1 vssd1 vccd1 vccd1 _18628_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09361_ _11484_/B1 _09352_/X _11466_/B1 vssd1 vssd1 vccd1 vccd1 _09361_/X sky130_fd_sc_hd__a21o_1
XFILLER_212_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18559_ _19613_/CLK _18559_/D vssd1 vssd1 vccd1 vccd1 _18559_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19134_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09292_ _12389_/A1 _09290_/X _09291_/X vssd1 vssd1 vccd1 vccd1 _09292_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _14837_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _15000_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 _09002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 _09401_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_56 _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_67 _10238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_89 _10459_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09628_ _18599_/Q _18170_/Q _10313_/S vssd1 vssd1 vccd1 vccd1 _09628_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09559_ _17914_/Q _09643_/A _09558_/Y _09367_/B vssd1 vssd1 vccd1 vccd1 _09561_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _12570_/A _12570_/B _12570_/C _12570_/D vssd1 vssd1 vccd1 vccd1 _12570_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ _12625_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _13316_/A sky130_fd_sc_hd__and2_2
XFILLER_184_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11452_ _11452_/A _11452_/B vssd1 vssd1 vccd1 vccd1 _11452_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14240_ _18118_/Q _14244_/B vssd1 vssd1 vccd1 vccd1 _14240_/X sky130_fd_sc_hd__or2_1
XFILLER_109_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10403_ _10401_/X _10402_/X _10403_/S vssd1 vssd1 vccd1 vccd1 _10403_/X sky130_fd_sc_hd__mux2_1
X_14171_ _16892_/A _14171_/B vssd1 vssd1 vccd1 vccd1 _18083_/D sky130_fd_sc_hd__and2_1
X_11383_ _11459_/A1 _11381_/X _11382_/X _11459_/B1 vssd1 vssd1 vccd1 vccd1 _11383_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_165_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10334_ _10334_/A1 _19158_/Q _09179_/B _19126_/Q vssd1 vssd1 vccd1 vccd1 _10334_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13122_ _13122_/A vssd1 vssd1 vccd1 vccd1 _13122_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17930_ _17930_/CLK _17930_/D vssd1 vssd1 vccd1 vccd1 _17930_/Q sky130_fd_sc_hd__dfxtp_4
X_13053_ _13100_/A _13053_/B vssd1 vssd1 vccd1 vccd1 _17925_/D sky130_fd_sc_hd__and2_1
XFILLER_279_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10265_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10265_/X sky130_fd_sc_hd__or2_1
XFILLER_79_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12004_ _17771_/Q _17672_/A0 _12021_/S vssd1 vssd1 vccd1 vccd1 _17771_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1300 _12786_/X vssd1 vssd1 vccd1 vccd1 _12788_/B sky130_fd_sc_hd__buf_6
Xfanout1311 _11741_/A2 vssd1 vssd1 vccd1 vccd1 _14522_/A2 sky130_fd_sc_hd__clkbuf_4
X_17861_ _19273_/CLK _17861_/D vssd1 vssd1 vccd1 vccd1 _17861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1322 _10996_/B1 vssd1 vssd1 vccd1 vccd1 _11459_/B1 sky130_fd_sc_hd__clkbuf_16
X_10196_ _11411_/A _10196_/B vssd1 vssd1 vccd1 vccd1 _10196_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1333 _10265_/A vssd1 vssd1 vccd1 vccd1 _09683_/A sky130_fd_sc_hd__buf_6
Xfanout1344 _09853_/S vssd1 vssd1 vccd1 vccd1 _11084_/S sky130_fd_sc_hd__buf_8
X_16812_ _19293_/Q _16815_/C _16812_/B1 vssd1 vssd1 vccd1 vccd1 _16812_/Y sky130_fd_sc_hd__o21ai_1
Xfanout1355 _10841_/C1 vssd1 vssd1 vccd1 vccd1 _09919_/C1 sky130_fd_sc_hd__clkbuf_16
X_19600_ _19600_/CLK _19600_/D vssd1 vssd1 vccd1 vccd1 _19600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_282_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1366 _11309_/S vssd1 vssd1 vccd1 vccd1 _10940_/S sky130_fd_sc_hd__buf_4
XFILLER_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17792_ _19650_/CLK _17792_/D vssd1 vssd1 vccd1 vccd1 _17792_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_93_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1377 _11073_/B1 vssd1 vssd1 vccd1 vccd1 _09770_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_266_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1388 _09843_/S vssd1 vssd1 vccd1 vccd1 _11147_/S sky130_fd_sc_hd__buf_6
Xfanout1399 fanout1407/X vssd1 vssd1 vccd1 vccd1 _09671_/S sky130_fd_sc_hd__buf_6
X_19531_ _19531_/CLK _19531_/D vssd1 vssd1 vccd1 vccd1 _19531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_282_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16743_ _19267_/Q _19266_/Q _16743_/C vssd1 vssd1 vccd1 vccd1 _16746_/B sky130_fd_sc_hd__and3_1
X_13955_ _13637_/A _14036_/B _13941_/X vssd1 vssd1 vccd1 vccd1 _13955_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19462_ _19534_/CLK _19462_/D vssd1 vssd1 vccd1 vccd1 _19462_/Q sky130_fd_sc_hd__dfxtp_2
X_12906_ _08897_/A _15151_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _12906_/X sky130_fd_sc_hd__mux2_1
X_16674_ _19246_/Q _19245_/Q _16674_/C vssd1 vssd1 vccd1 vccd1 _16675_/C sky130_fd_sc_hd__and3_1
X_13886_ _13876_/Y _13885_/Y _13920_/B2 _13875_/X vssd1 vssd1 vccd1 vccd1 _13886_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18413_ _18632_/CLK _18413_/D vssd1 vssd1 vccd1 vccd1 _18413_/Q sky130_fd_sc_hd__dfxtp_1
X_15625_ _15661_/B _15625_/B _15625_/C vssd1 vssd1 vccd1 vccd1 _15625_/Y sky130_fd_sc_hd__nand3_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12837_/A _12837_/B vssd1 vssd1 vccd1 vccd1 _12837_/X sky130_fd_sc_hd__or2_1
X_19393_ _19525_/CLK _19393_/D vssd1 vssd1 vccd1 vccd1 _19393_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _19622_/CLK _18344_/D vssd1 vssd1 vccd1 vccd1 _18344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _15482_/Y _15508_/X _15557_/C _15555_/Y _15530_/Y vssd1 vssd1 vccd1 vccd1
+ _15556_/X sky130_fd_sc_hd__o311a_4
XFILLER_188_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12768_ _12768_/A _12768_/B vssd1 vssd1 vccd1 vccd1 _12857_/S sky130_fd_sc_hd__or2_1
XFILLER_159_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14507_ _17709_/A0 _18357_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _18357_/D sky130_fd_sc_hd__mux2_1
X_11719_ _14696_/A _15835_/A _14417_/B vssd1 vssd1 vccd1 vccd1 _11719_/X sky130_fd_sc_hd__or3b_4
X_18275_ _18593_/CLK _18275_/D vssd1 vssd1 vccd1 vccd1 _18275_/Q sky130_fd_sc_hd__dfxtp_1
X_15487_ _15487_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _15489_/B sky130_fd_sc_hd__nor2_1
X_12699_ _12695_/X _12698_/X _12943_/S vssd1 vssd1 vccd1 vccd1 _12699_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17226_ _19426_/Q _17256_/B vssd1 vssd1 vccd1 vccd1 _17226_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput10 core_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_2
X_14438_ _18577_/Q _14451_/B vssd1 vssd1 vccd1 vccd1 _18290_/D sky130_fd_sc_hd__and2_1
Xinput21 core_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_2
Xinput32 core_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_2
Xinput43 dout0[0] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_2
XFILLER_128_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput54 dout0[1] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_2
X_17157_ _17157_/A _17583_/A vssd1 vssd1 vccd1 vccd1 _17453_/A sky130_fd_sc_hd__nand2_1
Xinput65 dout0[2] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_2
X_14369_ _18221_/Q _16543_/A0 _14383_/S vssd1 vssd1 vccd1 vccd1 _18221_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput76 dout0[3] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_2
Xinput87 dout0[4] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_2
X_16108_ _16142_/A1 _16107_/Y _16149_/A vssd1 vssd1 vccd1 vccd1 _18756_/D sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_137_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19304_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput98 dout0[5] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17088_ _17172_/B _17108_/A2 _17087_/X _17350_/A vssd1 vssd1 vccd1 vccd1 _19377_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08930_ _08914_/X _11985_/C _08927_/Y _08929_/X vssd1 vssd1 vccd1 vccd1 _08930_/Y
+ sky130_fd_sc_hd__a211oi_4
X_16039_ _16054_/A _18738_/Q _16063_/A vssd1 vssd1 vccd1 vccd1 _16039_/X sky130_fd_sc_hd__or3_2
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08861_ _16075_/A vssd1 vssd1 vccd1 vccd1 _08861_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09413_ _10294_/A1 _18140_/Q _18786_/Q _09428_/B2 vssd1 vssd1 vccd1 vccd1 _09413_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_280_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09344_ _18024_/Q _17992_/Q _09344_/S vssd1 vssd1 vccd1 vccd1 _09344_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09275_ _11484_/B1 _09266_/X _11466_/B1 vssd1 vssd1 vccd1 vccd1 _09275_/X sky130_fd_sc_hd__a21o_1
XFILLER_178_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _18626_/Q _10054_/S vssd1 vssd1 vccd1 vccd1 _10050_/X sky130_fd_sc_hd__or2_1
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13740_ _13938_/A _13740_/B vssd1 vssd1 vccd1 vccd1 _13740_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10952_ _11358_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _10952_/Y sky130_fd_sc_hd__nand2_1
XFILLER_232_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13671_ _13259_/X _13663_/X _13666_/Y _13670_/X vssd1 vssd1 vccd1 vccd1 _13671_/X
+ sky130_fd_sc_hd__a31o_1
X_10883_ _11594_/A1 _18959_/Q _18224_/Q _11613_/S vssd1 vssd1 vccd1 vccd1 _10883_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15410_ _15456_/C _15410_/B vssd1 vssd1 vccd1 vccd1 _15410_/Y sky130_fd_sc_hd__xnor2_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ _12622_/A _13226_/A vssd1 vssd1 vccd1 vccd1 _13261_/B sky130_fd_sc_hd__nand2_1
X_16390_ _16490_/A0 _19001_/Q _16390_/S vssd1 vssd1 vccd1 vccd1 _19001_/D sky130_fd_sc_hd__mux2_1
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15341_ _18573_/Q _15342_/B vssd1 vssd1 vccd1 vccd1 _15388_/C sky130_fd_sc_hd__and2_2
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12553_ _12553_/A _12553_/B _12553_/C _12553_/D vssd1 vssd1 vccd1 vccd1 _12563_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18060_ _19142_/CLK _18060_/D vssd1 vssd1 vccd1 vccd1 _18060_/Q sky130_fd_sc_hd__dfxtp_1
X_11504_ _11511_/A _11504_/B vssd1 vssd1 vccd1 vccd1 _11509_/A sky130_fd_sc_hd__and2_1
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15272_ _15314_/C _15272_/B vssd1 vssd1 vccd1 vccd1 _15272_/X sky130_fd_sc_hd__or2_1
XFILLER_185_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12484_ _12488_/A _17918_/Q _12483_/Y vssd1 vssd1 vccd1 vccd1 _12553_/B sky130_fd_sc_hd__a21o_2
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17011_ _19342_/Q _17043_/B vssd1 vssd1 vccd1 vccd1 _17011_/X sky130_fd_sc_hd__or2_1
XFILLER_172_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14223_ _18283_/Q _14261_/A2 _14222_/X _15718_/C1 vssd1 vssd1 vccd1 vccd1 _18109_/D
+ sky130_fd_sc_hd__o211a_1
X_11435_ _11512_/A1 _18607_/Q _18178_/Q _11513_/B2 vssd1 vssd1 vccd1 vccd1 _11435_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11366_ _09141_/A _15404_/A _11337_/X vssd1 vssd1 vccd1 vccd1 _12596_/B sky130_fd_sc_hd__o21ai_4
X_14154_ _14153_/B _14153_/C _14153_/D _14154_/B1 vssd1 vssd1 vccd1 vccd1 _14158_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13105_ _17830_/Q _13105_/B vssd1 vssd1 vccd1 vccd1 _13105_/Y sky130_fd_sc_hd__nor2_1
X_10317_ _10323_/A1 _19222_/Q _19190_/Q _10687_/S _11480_/C1 vssd1 vssd1 vccd1 vccd1
+ _10317_/X sky130_fd_sc_hd__a221o_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14085_ _16204_/A0 _18025_/Q _14106_/S vssd1 vssd1 vccd1 vccd1 _18025_/D sky130_fd_sc_hd__mux2_1
X_11297_ _09050_/X _09489_/B _11296_/Y _09030_/X vssd1 vssd1 vccd1 vccd1 _11297_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18962_ _19154_/CLK _18962_/D vssd1 vssd1 vccd1 vccd1 _18962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10248_ _18264_/Q _18839_/Q _10253_/C vssd1 vssd1 vccd1 vccd1 _10248_/X sky130_fd_sc_hd__mux2_1
X_17913_ _19206_/CLK _17913_/D vssd1 vssd1 vccd1 vccd1 _17913_/Q sky130_fd_sc_hd__dfxtp_4
X_13036_ _11740_/A _13349_/B _13035_/Y _13227_/C1 vssd1 vssd1 vccd1 vccd1 _13036_/X
+ sky130_fd_sc_hd__a211o_1
X_18893_ _19075_/CLK _18893_/D vssd1 vssd1 vccd1 vccd1 _18893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1130 _12322_/Y vssd1 vssd1 vccd1 vccd1 _15751_/A sky130_fd_sc_hd__buf_6
XFILLER_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1141 _11333_/A1 vssd1 vssd1 vccd1 vccd1 _10532_/A sky130_fd_sc_hd__buf_6
XFILLER_79_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17844_ _19470_/CLK _17844_/D vssd1 vssd1 vccd1 vccd1 _17844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_266_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10179_ _10169_/X _10172_/X _10175_/X _10178_/X _10243_/A _09264_/S vssd1 vssd1 vccd1
+ vccd1 _10180_/B sky130_fd_sc_hd__mux4_2
Xfanout1152 _13622_/A vssd1 vssd1 vccd1 vccd1 _13254_/B2 sky130_fd_sc_hd__buf_2
Xfanout1163 _15852_/X vssd1 vssd1 vccd1 vccd1 _15908_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1174 _15850_/X vssd1 vssd1 vccd1 vccd1 _15946_/A2 sky130_fd_sc_hd__buf_2
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1185 _15303_/B vssd1 vssd1 vccd1 vccd1 _15426_/B sky130_fd_sc_hd__buf_6
XFILLER_120_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1196 _16877_/B1 vssd1 vssd1 vccd1 vccd1 _16893_/B1 sky130_fd_sc_hd__buf_2
X_17775_ _18613_/CLK _17775_/D vssd1 vssd1 vccd1 vccd1 _17775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14987_ input64/X input100/X _15007_/S vssd1 vssd1 vccd1 vccd1 _14988_/A sky130_fd_sc_hd__mux2_2
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16726_ _19261_/Q _16728_/C _16725_/Y vssd1 vssd1 vccd1 vccd1 _19261_/D sky130_fd_sc_hd__o21a_1
X_19514_ _19546_/CLK _19514_/D vssd1 vssd1 vccd1 vccd1 _19514_/Q sky130_fd_sc_hd__dfxtp_1
X_13938_ _13938_/A _13938_/B vssd1 vssd1 vccd1 vccd1 _13938_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19445_ _19531_/CLK _19445_/D vssd1 vssd1 vccd1 vccd1 _19445_/Q sky130_fd_sc_hd__dfxtp_2
X_16657_ _19241_/Q _16661_/C vssd1 vssd1 vccd1 vccd1 _16659_/B sky130_fd_sc_hd__nor2_1
X_13869_ _15133_/A _13867_/X _13868_/Y _13869_/B2 vssd1 vssd1 vccd1 vccd1 _13870_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_234_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15608_ _19478_/Q _19412_/Q vssd1 vssd1 vccd1 vccd1 _15610_/A sky130_fd_sc_hd__and2_1
XFILLER_210_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19376_ _19543_/CLK _19376_/D vssd1 vssd1 vccd1 vccd1 _19376_/Q sky130_fd_sc_hd__dfxtp_1
X_16588_ _16621_/A0 _19192_/Q _16589_/S vssd1 vssd1 vccd1 vccd1 _19192_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18327_ _19649_/CLK _18327_/D vssd1 vssd1 vccd1 vccd1 _18327_/Q sky130_fd_sc_hd__dfxtp_1
X_15539_ _19443_/Q _15661_/B _17199_/A vssd1 vssd1 vccd1 vccd1 _15539_/X sky130_fd_sc_hd__o21a_1
XFILLER_176_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ _17900_/Q _12442_/B vssd1 vssd1 vccd1 vccd1 _12264_/B sky130_fd_sc_hd__nand2_8
X_18258_ _19025_/CLK _18258_/D vssd1 vssd1 vccd1 vccd1 _18258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ _19421_/Q fanout533/X _17208_/Y _17119_/B vssd1 vssd1 vccd1 vccd1 _17210_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_163_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18189_ _19641_/CLK _18189_/D vssd1 vssd1 vccd1 vccd1 _18189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09962_ _09960_/X _09961_/X _10300_/S vssd1 vssd1 vccd1 vccd1 _09962_/X sky130_fd_sc_hd__mux2_1
X_08913_ _14741_/A _08907_/Y _08912_/Y _08991_/A vssd1 vssd1 vccd1 vccd1 _08913_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _11286_/B1 _09877_/Y _09892_/X vssd1 vssd1 vccd1 vccd1 _09893_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_281_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08844_ _10253_/A vssd1 vssd1 vccd1 vccd1 _08844_/Y sky130_fd_sc_hd__inv_2
XFILLER_273_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19201_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_508 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_519 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09327_ _09027_/A _10085_/B _09322_/X _09030_/X vssd1 vssd1 vccd1 vccd1 _09327_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_240_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09258_ _18025_/Q _17993_/Q _09269_/S vssd1 vssd1 vccd1 vccd1 _09258_/X sky130_fd_sc_hd__mux2_1
XFILLER_279_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09189_ _11332_/B1 _09188_/X _11257_/C1 vssd1 vssd1 vccd1 vccd1 _09189_/X sky130_fd_sc_hd__o21a_1
XFILLER_135_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11220_ _09019_/Y _10605_/X _09030_/X vssd1 vssd1 vccd1 vccd1 _11220_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ _09683_/A _11149_/X _11150_/X _09106_/B vssd1 vssd1 vccd1 vccd1 _11151_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10102_ _18873_/Q _10176_/S _10101_/X _11397_/A1 vssd1 vssd1 vccd1 vccd1 _10102_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ _18456_/Q _18357_/Q _11309_/S vssd1 vssd1 vccd1 vccd1 _11082_/X sky130_fd_sc_hd__mux2_1
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput200 localMemory_wb_adr_i[19] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput211 localMemory_wb_adr_i[7] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14910_ _18492_/Q _15011_/A2 _14909_/Y _16803_/A vssd1 vssd1 vccd1 vccd1 _18492_/D
+ sky130_fd_sc_hd__a211o_1
Xinput222 localMemory_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input222/X sky130_fd_sc_hd__buf_8
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10033_ _10031_/X _10032_/X _10033_/S vssd1 vssd1 vccd1 vccd1 _10033_/X sky130_fd_sc_hd__mux2_1
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput233 localMemory_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 input233/X sky130_fd_sc_hd__clkbuf_16
XFILLER_237_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15890_ _15890_/A _15905_/B _15905_/C vssd1 vssd1 vccd1 vccd1 _15890_/X sky130_fd_sc_hd__and3_1
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput244 localMemory_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input244/X sky130_fd_sc_hd__buf_8
Xinput255 manufacturerID[1] vssd1 vssd1 vccd1 vccd1 _15860_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput266 partID[11] vssd1 vssd1 vccd1 vccd1 _15923_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput277 partID[7] vssd1 vssd1 vccd1 vccd1 _15911_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14841_ _14839_/X _14840_/X _14714_/B vssd1 vssd1 vccd1 vccd1 _14841_/X sky130_fd_sc_hd__a21o_1
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _17117_/B _17589_/B _17558_/X _17603_/B1 vssd1 vssd1 vccd1 vccd1 _19522_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ _18109_/Q _14801_/B _14770_/X _14771_/X vssd1 vssd1 vccd1 vccd1 _14772_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_263_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11984_ _18738_/Q _18730_/Q _16056_/B _15849_/A _11983_/X vssd1 vssd1 vccd1 vccd1
+ _11984_/X sky130_fd_sc_hd__a32o_4
XFILLER_44_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16511_ _17644_/A0 _19117_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _19117_/D sky130_fd_sc_hd__mux2_1
XFILLER_217_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13723_ _13713_/Y _13722_/Y _13747_/B2 _13712_/X vssd1 vssd1 vccd1 vccd1 _13723_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_260_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10935_ _11328_/S _10930_/X _10934_/X _11579_/A vssd1 vssd1 vccd1 vccd1 _10935_/X
+ sky130_fd_sc_hd__o211a_1
X_17491_ _18582_/Q _17544_/A _08883_/A vssd1 vssd1 vccd1 vccd1 _17491_/X sky130_fd_sc_hd__o21a_1
XFILLER_210_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19230_ _19319_/CLK _19230_/D vssd1 vssd1 vccd1 vccd1 _19230_/Q sky130_fd_sc_hd__dfxtp_4
X_16442_ _19050_/Q _16607_/A0 _16458_/S vssd1 vssd1 vccd1 vccd1 _19050_/D sky130_fd_sc_hd__mux2_1
X_13654_ _19414_/Q _13654_/A2 _13654_/B1 vssd1 vssd1 vccd1 vccd1 _13654_/X sky130_fd_sc_hd__a21o_1
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10866_ _10864_/X _10865_/X _10866_/S vssd1 vssd1 vccd1 vccd1 _10866_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19161_ _19628_/CLK _19161_/D vssd1 vssd1 vccd1 vccd1 _19161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _09984_/A _09984_/B _12842_/A _12842_/B vssd1 vssd1 vccd1 vccd1 _12900_/B
+ sky130_fd_sc_hd__a22oi_4
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _17705_/A0 _18984_/Q _16390_/S vssd1 vssd1 vccd1 vccd1 _18984_/D sky130_fd_sc_hd__mux2_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _17875_/Q _13747_/A2 _13584_/X _13682_/B2 vssd1 vssd1 vccd1 vccd1 _13585_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10797_ _10795_/X _10796_/X _11358_/A vssd1 vssd1 vccd1 vccd1 _10797_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _19450_/CLK _18112_/D vssd1 vssd1 vccd1 vccd1 _18112_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15324_ _15324_/A _15324_/B vssd1 vssd1 vccd1 vccd1 _15324_/X sky130_fd_sc_hd__xor2_1
X_12536_ _12579_/A _12552_/B vssd1 vssd1 vccd1 vccd1 _12536_/Y sky130_fd_sc_hd__nor2_8
X_19092_ _19092_/CLK _19092_/D vssd1 vssd1 vccd1 vccd1 _19092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18043_ _19613_/CLK _18043_/D vssd1 vssd1 vccd1 vccd1 _18043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15255_ _19463_/Q _15254_/Y _15400_/S vssd1 vssd1 vccd1 vccd1 _15255_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12467_ _12499_/A _12513_/B vssd1 vssd1 vccd1 vccd1 _12507_/A sky130_fd_sc_hd__nor2_4
XFILLER_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14206_ _18101_/Q _14266_/B vssd1 vssd1 vccd1 vccd1 _14206_/X sky130_fd_sc_hd__or2_1
X_11418_ _11511_/A _11413_/X _11417_/X vssd1 vssd1 vccd1 vccd1 _11418_/Y sky130_fd_sc_hd__a21oi_2
X_15186_ _19460_/Q _19394_/Q vssd1 vssd1 vccd1 vccd1 _15186_/Y sky130_fd_sc_hd__nor2_1
X_12398_ _12962_/A0 _12427_/A _12397_/Y _12428_/C1 vssd1 vssd1 vccd1 vccd1 _17907_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14137_ _16488_/A0 _18076_/Q _14137_/S vssd1 vssd1 vccd1 vccd1 _18076_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11349_ _11606_/S _11346_/X _11348_/X vssd1 vssd1 vccd1 vccd1 _11349_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_98_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14068_ _17685_/A0 _18010_/Q _14072_/S vssd1 vssd1 vccd1 vccd1 _18010_/D sky130_fd_sc_hd__mux2_1
X_18945_ _19147_/CLK _18945_/D vssd1 vssd1 vccd1 vccd1 _18945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13019_ _19365_/Q _13247_/A2 _13017_/X _13018_/X _13247_/C1 vssd1 vssd1 vccd1 vccd1
+ _13019_/X sky130_fd_sc_hd__o221a_4
XFILLER_140_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18876_ _19619_/CLK _18876_/D vssd1 vssd1 vccd1 vccd1 _18876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17827_ _18713_/CLK _17827_/D vssd1 vssd1 vccd1 vccd1 _17827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17758_ _19586_/CLK _17758_/D vssd1 vssd1 vccd1 vccd1 _17758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16709_ _19255_/Q _16706_/B _16707_/Y vssd1 vssd1 vccd1 vccd1 _19255_/D sky130_fd_sc_hd__o21a_1
X_17689_ _17722_/A0 _19616_/Q _17689_/S vssd1 vssd1 vccd1 vccd1 _19616_/D sky130_fd_sc_hd__mux2_1
XFILLER_207_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19428_ _19492_/CLK _19428_/D vssd1 vssd1 vccd1 vccd1 _19428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19359_ _19540_/CLK _19359_/D vssd1 vssd1 vccd1 vccd1 _19359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09112_ _09109_/X _09111_/X _12408_/A vssd1 vssd1 vccd1 vccd1 _09112_/X sky130_fd_sc_hd__a21bo_1
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_152_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19466_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_164_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09043_ _09043_/A _11217_/A _11217_/B vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__and3_4
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout901 _16204_/A0 vssd1 vssd1 vccd1 vccd1 _17668_/A0 sky130_fd_sc_hd__buf_2
XFILLER_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09945_ _10471_/S _10027_/B vssd1 vssd1 vccd1 vccd1 _09945_/Y sky130_fd_sc_hd__nand2_1
Xfanout912 _16385_/S vssd1 vssd1 vccd1 vccd1 _16391_/S sky130_fd_sc_hd__buf_8
Xfanout923 _16227_/Y vssd1 vssd1 vccd1 vccd1 _16245_/S sky130_fd_sc_hd__buf_8
Xfanout934 _14983_/B1 vssd1 vssd1 vccd1 vccd1 _14973_/B1 sky130_fd_sc_hd__buf_4
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout945 _14670_/Y vssd1 vssd1 vccd1 vccd1 _14714_/B sky130_fd_sc_hd__buf_4
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout956 _14599_/X vssd1 vssd1 vccd1 vccd1 _14628_/S sky130_fd_sc_hd__buf_12
Xfanout967 _14104_/S vssd1 vssd1 vccd1 vccd1 _14106_/S sky130_fd_sc_hd__buf_12
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09876_ _10030_/C1 _09872_/X _09875_/X vssd1 vssd1 vccd1 vccd1 _09877_/B sky130_fd_sc_hd__a21oi_1
XFILLER_246_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout978 _13115_/B2 vssd1 vssd1 vccd1 vccd1 _13945_/B2 sky130_fd_sc_hd__buf_6
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _16034_/S vssd1 vssd1 vccd1 vccd1 _16069_/A sky130_fd_sc_hd__inv_2
XFILLER_58_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_305 _18113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_316 _18125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_327 _11957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 _11482_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_349 _15481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ _11277_/A1 _19576_/Q _10370_/S _19608_/Q _10371_/S vssd1 vssd1 vccd1 vccd1
+ _10720_/X sky130_fd_sc_hd__o221a_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10651_ _10662_/A1 _18227_/Q _10650_/S _18962_/Q _10668_/S vssd1 vssd1 vccd1 vccd1
+ _10651_/X sky130_fd_sc_hd__o221a_1
XFILLER_179_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _17837_/Q _13844_/A2 _13844_/B1 _17869_/Q vssd1 vssd1 vccd1 vccd1 _13370_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10582_ _18618_/Q _18189_/Q _10582_/S vssd1 vssd1 vccd1 vccd1 _10582_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12321_ _17915_/Q _12321_/B _17917_/Q _17916_/Q vssd1 vssd1 vccd1 vccd1 _12323_/B
+ sky130_fd_sc_hd__or4bb_4
XFILLER_182_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15040_ _18529_/Q _17342_/A _11711_/A _11711_/B _16627_/S vssd1 vssd1 vccd1 vccd1
+ _18529_/D sky130_fd_sc_hd__a41o_1
X_12252_ _17883_/Q _12253_/C _12251_/Y vssd1 vssd1 vccd1 vccd1 _17883_/D sky130_fd_sc_hd__o21a_1
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11203_ _11618_/A1 _19602_/Q _19570_/Q _10726_/S vssd1 vssd1 vccd1 vccd1 _11203_/X
+ sky130_fd_sc_hd__a22o_1
X_12183_ _17857_/Q _12184_/C _17858_/Q vssd1 vssd1 vccd1 vccd1 _12185_/B sky130_fd_sc_hd__a21oi_1
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11134_ _15478_/A vssd1 vssd1 vccd1 vccd1 _11134_/Y sky130_fd_sc_hd__inv_2
X_16991_ _19332_/Q _17009_/B vssd1 vssd1 vccd1 vccd1 _16991_/X sky130_fd_sc_hd__or2_1
XFILLER_205_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15942_ _18689_/Q _15948_/A2 _15948_/B1 _15941_/X _15948_/C1 vssd1 vssd1 vccd1 vccd1
+ _15942_/X sky130_fd_sc_hd__a221o_1
X_11065_ _17969_/Q _11295_/A2 _11216_/B1 vssd1 vssd1 vccd1 vccd1 _11066_/B sky130_fd_sc_hd__a21oi_1
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18730_ _18738_/CLK _18730_/D vssd1 vssd1 vccd1 vccd1 _18730_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10016_ _11579_/A _10012_/X _10015_/X _10557_/S _11570_/B1 vssd1 vssd1 vccd1 vccd1
+ _10016_/X sky130_fd_sc_hd__o221a_1
X_18661_ _18666_/CLK _18661_/D vssd1 vssd1 vccd1 vccd1 _18661_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15873_ _18666_/Q _15853_/Y _15906_/B1 vssd1 vssd1 vccd1 vccd1 _15873_/X sky130_fd_sc_hd__a21o_1
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824_ input47/X input82/X _14844_/S vssd1 vssd1 vccd1 vccd1 _14825_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17612_ _19547_/Q _17624_/A2 _17591_/X _17196_/B _17611_/X vssd1 vssd1 vccd1 vccd1
+ _19547_/D sky130_fd_sc_hd__o221a_1
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _19453_/CLK _18592_/D vssd1 vssd1 vccd1 vccd1 _18592_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_221_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17543_ _13938_/B _17531_/B _17543_/B1 _17820_/Q vssd1 vssd1 vccd1 vccd1 _17544_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14755_ input103/X input74/X _14784_/S vssd1 vssd1 vccd1 vccd1 _14755_/X sky130_fd_sc_hd__mux2_8
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11967_ _18513_/Q _11720_/X _11917_/X _11968_/B2 vssd1 vssd1 vccd1 vccd1 _11967_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13706_ _13736_/B _13706_/B vssd1 vssd1 vccd1 vccd1 _13706_/X sky130_fd_sc_hd__or2_1
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17474_ _19506_/Q _17547_/B _17472_/X _17473_/Y _17350_/A vssd1 vssd1 vccd1 vccd1
+ _19506_/D sky130_fd_sc_hd__o221a_1
X_10918_ _11305_/A1 _18223_/Q _11094_/S _18958_/Q _10918_/C1 vssd1 vssd1 vccd1 vccd1
+ _10918_/X sky130_fd_sc_hd__o221a_1
XFILLER_189_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14686_ _19227_/Q _14934_/C vssd1 vssd1 vccd1 vccd1 _15834_/B sky130_fd_sc_hd__nand2_4
XFILLER_204_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11898_ _11826_/B _11875_/Y _11897_/X vssd1 vssd1 vccd1 vccd1 _11899_/C sky130_fd_sc_hd__o21ai_2
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19213_ _19213_/CLK _19213_/D vssd1 vssd1 vccd1 vccd1 _19213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16425_ _17723_/A0 _19034_/Q _16425_/S vssd1 vssd1 vccd1 vccd1 _19034_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13637_ _13637_/A _14016_/B vssd1 vssd1 vccd1 vccd1 _13637_/X sky130_fd_sc_hd__or2_4
X_10849_ _10850_/A1 _19574_/Q _10853_/S _19606_/Q _11311_/C1 vssd1 vssd1 vccd1 vccd1
+ _10849_/X sky130_fd_sc_hd__o221a_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19144_ _19630_/CLK _19144_/D vssd1 vssd1 vccd1 vccd1 _19144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16356_ _18968_/Q _17688_/A0 _16357_/S vssd1 vssd1 vccd1 vccd1 _18968_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13568_ _13568_/A _13568_/B vssd1 vssd1 vccd1 vccd1 _14148_/A sky130_fd_sc_hd__xnor2_2
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15307_ _15307_/A _15307_/B _15305_/X vssd1 vssd1 vccd1 vccd1 _15308_/B sky130_fd_sc_hd__or3b_4
X_19075_ _19075_/CLK _19075_/D vssd1 vssd1 vccd1 vccd1 _19075_/Q sky130_fd_sc_hd__dfxtp_1
X_12519_ _12584_/A _12577_/B vssd1 vssd1 vccd1 vccd1 _12771_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16287_ _17718_/A0 _18901_/Q _16292_/S vssd1 vssd1 vccd1 vccd1 _18901_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13499_ _19409_/Q _13654_/A2 _13654_/B1 vssd1 vssd1 vccd1 vccd1 _13499_/X sky130_fd_sc_hd__a21o_1
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18026_ _19564_/CLK _18026_/D vssd1 vssd1 vccd1 vccd1 _18026_/Q sky130_fd_sc_hd__dfxtp_1
X_15238_ _15238_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _15238_/X sky130_fd_sc_hd__and2_1
XFILLER_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _17219_/A _15168_/X _15163_/Y _15424_/C1 vssd1 vssd1 vccd1 vccd1 _15169_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_126_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09730_ _11495_/B1 _09728_/X _09729_/X _09715_/X vssd1 vssd1 vccd1 vccd1 _09730_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_274_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18928_ _19639_/CLK _18928_/D vssd1 vssd1 vccd1 vccd1 _18928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09661_ _11556_/C _09650_/X _09660_/X _11687_/A vssd1 vssd1 vccd1 vccd1 _09661_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_269_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18859_ _19634_/CLK _18859_/D vssd1 vssd1 vccd1 vccd1 _18859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09592_ _10747_/A1 _09591_/X _09587_/X _08903_/A vssd1 vssd1 vccd1 vccd1 _09608_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_131_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09026_ _11218_/A _09048_/A vssd1 vssd1 vccd1 vccd1 _10085_/B sky130_fd_sc_hd__nand2_4
XFILLER_136_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1707 _08843_/Y vssd1 vssd1 vccd1 vccd1 _09350_/S sky130_fd_sc_hd__buf_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1718 _08828_/Y vssd1 vssd1 vccd1 vccd1 _16898_/A1 sky130_fd_sc_hd__buf_4
Xfanout720 _12497_/Y vssd1 vssd1 vccd1 vccd1 _13744_/B1 sky130_fd_sc_hd__buf_4
XFILLER_172_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout731 _11451_/X vssd1 vssd1 vccd1 vccd1 _11452_/B sky130_fd_sc_hd__buf_4
Xfanout1729 _08828_/A vssd1 vssd1 vccd1 vccd1 _12483_/A sky130_fd_sc_hd__buf_6
XFILLER_277_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09928_ _09457_/B _18876_/Q _09285_/C _11481_/A vssd1 vssd1 vccd1 vccd1 _09928_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout742 _17641_/A0 vssd1 vssd1 vccd1 vccd1 _17674_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_213_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout753 _13390_/S vssd1 vssd1 vccd1 vccd1 _13315_/S sky130_fd_sc_hd__buf_6
XFILLER_213_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout764 _09054_/X vssd1 vssd1 vccd1 vccd1 _09105_/A sky130_fd_sc_hd__buf_4
XFILLER_219_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout775 _17654_/S vssd1 vssd1 vccd1 vccd1 _17656_/S sky130_fd_sc_hd__buf_12
Xfanout786 _16525_/Y vssd1 vssd1 vccd1 vccd1 _16548_/S sky130_fd_sc_hd__buf_6
XFILLER_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout797 _16325_/S vssd1 vssd1 vccd1 vccd1 _16320_/S sky130_fd_sc_hd__buf_12
X_09859_ _09859_/A _09859_/B _09859_/C vssd1 vssd1 vccd1 vccd1 _09859_/Y sky130_fd_sc_hd__nand3_4
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12870_ _13421_/A _11732_/Y _12761_/B _12869_/A _13185_/A vssd1 vssd1 vccd1 vccd1
+ _12870_/X sky130_fd_sc_hd__a221o_1
XFILLER_246_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _11819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _11807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ _11820_/A _11819_/X _11820_/Y _11859_/B vssd1 vssd1 vccd1 vccd1 _11822_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_124 _11825_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _11831_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _11868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _11904_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14596_/A _14540_/B vssd1 vssd1 vccd1 vccd1 _18378_/D sky130_fd_sc_hd__or2_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _18571_/Q _11759_/A2 _11844_/A _11751_/Y vssd1 vssd1 vccd1 vccd1 _11752_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _13988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_179 _13513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10703_ _11161_/S _10698_/X _10702_/X vssd1 vssd1 vccd1 vccd1 _10703_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14471_ _18323_/Q _17708_/A0 _14477_/S vssd1 vssd1 vccd1 vccd1 _18323_/D sky130_fd_sc_hd__mux2_1
XFILLER_202_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _13366_/B _11683_/B _11664_/B vssd1 vssd1 vccd1 vccd1 _11684_/D sky130_fd_sc_hd__or3b_1
X_16210_ _17707_/A0 _18826_/Q _16212_/S vssd1 vssd1 vccd1 vccd1 _18826_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13422_ _15426_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13438_/B sky130_fd_sc_hd__nand2_1
XFILLER_220_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17190_ _17202_/A _17190_/B vssd1 vssd1 vccd1 vccd1 _17508_/A sky130_fd_sc_hd__nand2_2
X_10634_ _18649_/Q _18071_/Q _19090_/Q _18994_/Q _10634_/S0 _10918_/C1 vssd1 vssd1
+ vccd1 vccd1 _10634_/X sky130_fd_sc_hd__mux4_1
XFILLER_197_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _18773_/Q _16141_/B vssd1 vssd1 vccd1 vccd1 _16141_/Y sky130_fd_sc_hd__nand2_1
X_13353_ _13390_/S _12889_/X _13413_/B1 vssd1 vssd1 vccd1 vccd1 _13353_/X sky130_fd_sc_hd__a21o_1
X_10565_ _11583_/A _11135_/S _11181_/B1 _10564_/Y vssd1 vssd1 vccd1 vccd1 _10602_/A
+ sky130_fd_sc_hd__o22a_4
X_12304_ _11715_/C _12305_/B1 _12303_/X _12276_/X vssd1 vssd1 vccd1 vccd1 _14687_/A
+ sky130_fd_sc_hd__a22o_2
X_16072_ _16075_/A _16075_/C _16071_/Y vssd1 vssd1 vccd1 vccd1 _16072_/Y sky130_fd_sc_hd__o21ai_1
X_13284_ _17866_/Q _13847_/A2 _13722_/B1 _13283_/X vssd1 vssd1 vccd1 vccd1 _13284_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10496_ _18651_/Q _10496_/B vssd1 vssd1 vccd1 vccd1 _10496_/X sky130_fd_sc_hd__or2_1
XFILLER_182_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15023_ _18512_/Q input212/X _15024_/S vssd1 vssd1 vccd1 vccd1 _18512_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12235_ _12241_/A _12240_/C vssd1 vssd1 vccd1 vccd1 _12235_/Y sky130_fd_sc_hd__nor2_1
XFILLER_216_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12166_ _17851_/Q _12168_/C _12165_/Y vssd1 vssd1 vccd1 vccd1 _17851_/D sky130_fd_sc_hd__o21a_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ _11117_/A _11117_/B vssd1 vssd1 vccd1 vccd1 _11117_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12097_ _17826_/Q _12100_/C vssd1 vssd1 vccd1 vccd1 _12098_/B sky130_fd_sc_hd__and2_1
X_16974_ _17051_/D _17052_/B _17052_/C vssd1 vssd1 vccd1 vccd1 _16975_/C sky130_fd_sc_hd__or3_1
XFILLER_49_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18713_ _18713_/CLK _18713_/D vssd1 vssd1 vccd1 vccd1 _18713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15925_ _18684_/Q _15943_/A2 _15924_/X _15946_/C1 vssd1 vssd1 vccd1 vccd1 _18684_/D
+ sky130_fd_sc_hd__o211a_1
X_11048_ _11512_/A1 _18325_/Q _17776_/Q _11426_/B2 vssd1 vssd1 vccd1 vccd1 _11048_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_265_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 coreIndex[7] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_6
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15856_ _18661_/Q _15949_/A2 _15855_/X _14205_/A vssd1 vssd1 vccd1 vccd1 _18661_/D
+ sky130_fd_sc_hd__o211a_1
X_18644_ _19142_/CLK _18644_/D vssd1 vssd1 vccd1 vccd1 _18644_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_225_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14807_ _14803_/Y _14806_/X _14950_/B1 vssd1 vssd1 vccd1 vccd1 _14807_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15787_ _15787_/A _15787_/B vssd1 vssd1 vccd1 vccd1 _15788_/B sky130_fd_sc_hd__xnor2_1
X_18575_ _19433_/CLK _18575_/D vssd1 vssd1 vccd1 vccd1 _18575_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12999_ _13230_/A1 _12836_/Y _12999_/S vssd1 vssd1 vccd1 vccd1 _12999_/X sky130_fd_sc_hd__mux2_2
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14738_ _14718_/A _14737_/X _14846_/B1 vssd1 vssd1 vccd1 vccd1 _14738_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17526_ _18589_/Q _17544_/A vssd1 vssd1 vccd1 vccd1 _17526_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17457_ _17457_/A _17462_/B vssd1 vssd1 vccd1 vccd1 _17457_/Y sky130_fd_sc_hd__nand2_1
XFILLER_232_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14669_ _14688_/A _14669_/B vssd1 vssd1 vccd1 vccd1 _14680_/C sky130_fd_sc_hd__or2_2
XFILLER_221_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16408_ _17706_/A0 _19017_/Q _16420_/S vssd1 vssd1 vccd1 vccd1 _19017_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17388_ _12460_/A _15140_/B _17386_/X _17387_/X _14430_/B vssd1 vssd1 vccd1 vccd1
+ _19489_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16339_ _18951_/Q _17671_/A0 _16357_/S vssd1 vssd1 vccd1 vccd1 _18951_/D sky130_fd_sc_hd__mux2_1
X_19127_ _19203_/CLK _19127_/D vssd1 vssd1 vccd1 vccd1 _19127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19058_ _19219_/CLK _19058_/D vssd1 vssd1 vccd1 vccd1 _19058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput301 _11917_/X vssd1 vssd1 vccd1 vccd1 addr1[7] sky130_fd_sc_hd__buf_4
XFILLER_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput312 _11760_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[16] sky130_fd_sc_hd__buf_4
X_18009_ _19092_/CLK _18009_/D vssd1 vssd1 vccd1 vccd1 _18009_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput323 _11770_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[26] sky130_fd_sc_hd__buf_4
Xoutput334 _11784_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[0] sky130_fd_sc_hd__buf_4
XFILLER_126_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput345 _11787_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[1] sky130_fd_sc_hd__buf_4
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput356 _11789_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[2] sky130_fd_sc_hd__buf_4
Xoutput367 _11775_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[1] sky130_fd_sc_hd__buf_4
XFILLER_273_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput378 _11931_/X vssd1 vssd1 vccd1 vccd1 din0[11] sky130_fd_sc_hd__buf_4
Xoutput389 _11941_/X vssd1 vssd1 vccd1 vccd1 din0[21] sky130_fd_sc_hd__buf_4
XFILLER_141_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09713_ _09711_/X _09712_/X _10371_/S vssd1 vssd1 vccd1 vccd1 _09713_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09644_ _17913_/Q _09643_/A _09643_/Y _09367_/B vssd1 vssd1 vccd1 vccd1 _09647_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09575_ _11556_/C _09564_/X _09574_/X _11687_/A vssd1 vssd1 vccd1 vccd1 _09575_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10350_ _18075_/Q _10364_/B _10349_/X _10346_/S vssd1 vssd1 vccd1 vccd1 _10350_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_192_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09009_ _11691_/B1 _12409_/A2 _09008_/X _09650_/B1 _18396_/Q vssd1 vssd1 vccd1 vccd1
+ _09009_/X sky130_fd_sc_hd__o32a_2
X_10281_ _19095_/Q _18999_/Q _10281_/S vssd1 vssd1 vccd1 vccd1 _10281_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12020_ _17787_/Q _17688_/A0 _12021_/S vssd1 vssd1 vccd1 vccd1 _17787_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1504 _08968_/S0 vssd1 vssd1 vccd1 vccd1 _09973_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_120_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1515 fanout1524/X vssd1 vssd1 vccd1 vccd1 _09966_/S sky130_fd_sc_hd__buf_6
XFILLER_120_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1526 _11112_/A vssd1 vssd1 vccd1 vccd1 _11358_/A sky130_fd_sc_hd__buf_6
Xfanout1537 _10653_/A1 vssd1 vssd1 vccd1 vccd1 _10346_/S sky130_fd_sc_hd__buf_6
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout550 _17202_/A vssd1 vssd1 vccd1 vccd1 _17199_/A sky130_fd_sc_hd__buf_6
Xfanout1548 _10033_/S vssd1 vssd1 vccd1 vccd1 _11616_/S sky130_fd_sc_hd__clkbuf_8
Xfanout1559 _09381_/S vssd1 vssd1 vccd1 vccd1 _09374_/S sky130_fd_sc_hd__buf_8
Xfanout561 _15112_/Y vssd1 vssd1 vccd1 vccd1 _15537_/B1 sky130_fd_sc_hd__buf_4
XFILLER_265_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout572 _15124_/C vssd1 vssd1 vccd1 vccd1 _15381_/A3 sky130_fd_sc_hd__buf_6
XFILLER_120_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout583 _12338_/Y vssd1 vssd1 vccd1 vccd1 _12427_/A sky130_fd_sc_hd__buf_4
X_13971_ _15549_/A _13971_/A2 _13579_/A vssd1 vssd1 vccd1 vccd1 _13971_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout594 _14252_/B vssd1 vssd1 vccd1 vccd1 _14247_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_262_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15710_ _19451_/Q _15661_/B _17202_/A vssd1 vssd1 vccd1 vccd1 _15710_/X sky130_fd_sc_hd__o21a_1
XFILLER_247_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12922_ _13980_/B vssd1 vssd1 vccd1 vccd1 _12922_/Y sky130_fd_sc_hd__inv_2
X_16690_ _19249_/Q _19248_/Q _16690_/C _16690_/D vssd1 vssd1 vccd1 vccd1 _16699_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_246_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15641_ _15702_/A _15553_/B _15556_/X _15638_/X _15640_/Y vssd1 vssd1 vccd1 vccd1
+ _15641_/X sky130_fd_sc_hd__o221a_1
XFILLER_92_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12853_ _19394_/Q _12579_/Y _12771_/X _12852_/X _12581_/Y vssd1 vssd1 vccd1 vccd1
+ _12853_/X sky130_fd_sc_hd__a221o_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _19575_/CLK _18360_/D vssd1 vssd1 vccd1 vccd1 _18360_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11804_ _11804_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11804_/X sky130_fd_sc_hd__or2_4
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15572_ _15782_/A1 _15571_/X _15782_/B1 vssd1 vssd1 vccd1 vccd1 _15572_/X sky130_fd_sc_hd__a21o_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _13757_/A _13976_/B _12766_/X vssd1 vssd1 vccd1 vccd1 _12784_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_215_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _18131_/Q _17219_/A _17547_/A _17310_/B vssd1 vssd1 vccd1 vccd1 _17311_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _18406_/Q _14522_/Y _18372_/Q vssd1 vssd1 vccd1 vccd1 _14525_/B sky130_fd_sc_hd__o21ba_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18291_ _18593_/CLK _18291_/D vssd1 vssd1 vccd1 vccd1 _18291_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11735_/A _12957_/A vssd1 vssd1 vccd1 vccd1 _12956_/A sky130_fd_sc_hd__xnor2_4
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _14220_/A _17151_/A _17428_/A _17241_/B vssd1 vssd1 vccd1 vccd1 _17242_/X
+ sky130_fd_sc_hd__o22a_1
X_14454_ _14599_/A _16326_/A vssd1 vssd1 vccd1 vccd1 _14454_/Y sky130_fd_sc_hd__nor2_8
XFILLER_202_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11666_ _11666_/A _11727_/B vssd1 vssd1 vccd1 vccd1 _14347_/B sky130_fd_sc_hd__nor2_2
XFILLER_174_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13405_ _18116_/Q _13406_/B vssd1 vssd1 vccd1 vccd1 _13479_/C sky130_fd_sc_hd__and2_2
X_10617_ _18617_/Q _18188_/Q _10619_/S vssd1 vssd1 vccd1 vccd1 _10617_/X sky130_fd_sc_hd__mux2_1
X_17173_ _19409_/Q fanout534/X _17478_/A _17212_/B2 vssd1 vssd1 vccd1 vccd1 _17174_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14385_ _17692_/A0 _18236_/Q _14402_/S vssd1 vssd1 vccd1 vccd1 _18236_/D sky130_fd_sc_hd__mux2_1
XFILLER_259_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11597_ _18267_/Q _18842_/Q _11598_/S vssd1 vssd1 vccd1 vccd1 _11597_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16124_ _16140_/A1 _16123_/Y _16128_/B1 vssd1 vssd1 vccd1 vccd1 _18764_/D sky130_fd_sc_hd__a21oi_1
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13336_ _19535_/Q _19503_/Q _13372_/S vssd1 vssd1 vccd1 vccd1 _13336_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10548_ _11583_/A _10543_/X _10545_/X _10547_/X _11588_/B1 vssd1 vssd1 vccd1 vccd1
+ _10548_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16055_ _16055_/A vssd1 vssd1 vccd1 vccd1 _16063_/C sky130_fd_sc_hd__inv_2
X_13267_ _13267_/A _13316_/B vssd1 vssd1 vccd1 vccd1 _13267_/Y sky130_fd_sc_hd__nand2_1
X_10479_ _09853_/S _10474_/X _10478_/X vssd1 vssd1 vccd1 vccd1 _10479_/X sky130_fd_sc_hd__o21a_1
XFILLER_142_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15006_ _15006_/A1 _15005_/X _15006_/B1 vssd1 vssd1 vccd1 vccd1 _15006_/Y sky130_fd_sc_hd__o21ai_2
X_12218_ _17871_/Q _12218_/B vssd1 vssd1 vccd1 vccd1 _12224_/C sky130_fd_sc_hd__and2_2
XFILLER_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13198_ _13896_/B2 _13194_/X _13197_/X _12733_/S _13196_/Y vssd1 vssd1 vccd1 vccd1
+ _13198_/X sky130_fd_sc_hd__o221a_4
XFILLER_285_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12149_ _17845_/Q _12152_/C _17159_/A vssd1 vssd1 vccd1 vccd1 _12149_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_284_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16957_ _18770_/Q _16965_/A2 _16965_/B1 input235/X _16965_/C1 vssd1 vssd1 vccd1 vccd1
+ _16957_/X sky130_fd_sc_hd__a221o_1
XFILLER_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15908_ _15908_/A _15941_/S _15908_/C vssd1 vssd1 vccd1 vccd1 _15908_/X sky130_fd_sc_hd__and3_1
X_16888_ _16972_/A _16888_/B vssd1 vssd1 vccd1 vccd1 _19306_/D sky130_fd_sc_hd__and2_1
X_18627_ _18627_/CLK _18627_/D vssd1 vssd1 vccd1 vccd1 _18627_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15839_ _18743_/Q _12276_/A _16877_/B1 input226/X vssd1 vssd1 vccd1 vccd1 _15840_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_253_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09360_ _09360_/A _09360_/B vssd1 vssd1 vccd1 vccd1 _09360_/X sky130_fd_sc_hd__and2_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18558_ _19565_/CLK _18558_/D vssd1 vssd1 vccd1 vccd1 _18558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17509_ _19513_/Q _17523_/B _17507_/X _17508_/Y _17368_/A vssd1 vssd1 vccd1 vccd1
+ _19513_/D sky130_fd_sc_hd__o221a_1
X_09291_ _11498_/A1 _19204_/Q _19172_/Q _09290_/S _10144_/B1 vssd1 vssd1 vccd1 vccd1
+ _09291_/X sky130_fd_sc_hd__a221o_1
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18489_ _19286_/CLK _18489_/D vssd1 vssd1 vccd1 vccd1 _18489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 _14847_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_24 _15853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_35 _09002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_46 _09401_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19564_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_57 _12602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_68 _13843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09627_ _18241_/Q _18816_/Q _10313_/S vssd1 vssd1 vccd1 vccd1 _09627_/X sky130_fd_sc_hd__mux2_1
XFILLER_244_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09558_ _09643_/A _11798_/B vssd1 vssd1 vccd1 vccd1 _09558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09489_ _09574_/A _09489_/B _09489_/C vssd1 vssd1 vccd1 vccd1 _09489_/X sky130_fd_sc_hd__or3_2
XFILLER_168_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ _12625_/B vssd1 vssd1 vccd1 vccd1 _11522_/B sky130_fd_sc_hd__clkinv_2
XFILLER_157_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11451_ _17932_/Q _11451_/A2 _11450_/X _11451_/B2 vssd1 vssd1 vccd1 vccd1 _11451_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_183_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10402_ _11458_/A1 _17784_/Q _11462_/S _18333_/Q vssd1 vssd1 vccd1 vccd1 _10402_/X
+ sky130_fd_sc_hd__o22a_1
X_14170_ _18696_/Q _18083_/Q _14186_/S vssd1 vssd1 vccd1 vccd1 _14171_/B sky130_fd_sc_hd__mux2_1
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11382_ _11465_/A1 _19144_/Q _11384_/B _19112_/Q _10403_/S vssd1 vssd1 vccd1 vccd1
+ _11382_/X sky130_fd_sc_hd__o221a_1
X_13121_ _18108_/Q _13159_/C vssd1 vssd1 vccd1 vccd1 _13122_/A sky130_fd_sc_hd__xnor2_1
X_10333_ _10334_/A1 _18231_/Q _09179_/B _18966_/Q vssd1 vssd1 vccd1 vccd1 _10333_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13052_ _09562_/X _13292_/A2 _13051_/X _13256_/B1 _17925_/Q vssd1 vssd1 vccd1 vccd1
+ _13053_/B sky130_fd_sc_hd__a32o_1
X_10264_ _10262_/X _10263_/X _10264_/S vssd1 vssd1 vccd1 vccd1 _10265_/B sky130_fd_sc_hd__mux2_1
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12003_ _17770_/Q _17671_/A0 _12019_/S vssd1 vssd1 vccd1 vccd1 _17770_/D sky130_fd_sc_hd__mux2_1
XFILLER_278_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1301 _16969_/A2 vssd1 vssd1 vccd1 vccd1 _16965_/A2 sky130_fd_sc_hd__buf_4
XFILLER_279_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17860_ _18691_/CLK _17860_/D vssd1 vssd1 vccd1 vccd1 _17860_/Q sky130_fd_sc_hd__dfxtp_2
X_10195_ _11452_/A _10166_/X _10194_/Y _11023_/B1 vssd1 vssd1 vccd1 vccd1 _10196_/B
+ sky130_fd_sc_hd__o211ai_4
Xfanout1312 _11724_/Y vssd1 vssd1 vccd1 vccd1 _11741_/A2 sky130_fd_sc_hd__buf_4
Xfanout1323 _09099_/Y vssd1 vssd1 vccd1 vccd1 _10996_/B1 sky130_fd_sc_hd__buf_8
Xfanout1334 _10004_/A1 vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__buf_6
XFILLER_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16811_ _16811_/A _16811_/B _16815_/C vssd1 vssd1 vccd1 vccd1 _19292_/D sky130_fd_sc_hd__nor3_1
Xfanout1345 _09853_/S vssd1 vssd1 vccd1 vccd1 _11248_/S sky130_fd_sc_hd__buf_4
Xfanout1356 _09095_/Y vssd1 vssd1 vccd1 vccd1 _10841_/C1 sky130_fd_sc_hd__buf_6
XFILLER_282_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17791_ _19650_/CLK _17791_/D vssd1 vssd1 vccd1 vccd1 _17791_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1367 _10929_/S vssd1 vssd1 vccd1 vccd1 _11309_/S sky130_fd_sc_hd__clkbuf_8
Xfanout1378 _11073_/B1 vssd1 vssd1 vccd1 vccd1 _11094_/S sky130_fd_sc_hd__clkbuf_8
Xfanout1389 _09843_/S vssd1 vssd1 vccd1 vccd1 _10840_/S sky130_fd_sc_hd__buf_6
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19530_ _19530_/CLK _19530_/D vssd1 vssd1 vccd1 vccd1 _19530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16742_ _19267_/Q _16742_/B vssd1 vssd1 vccd1 vccd1 _16744_/B sky130_fd_sc_hd__nor2_1
XFILLER_207_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13954_ _14036_/B vssd1 vssd1 vccd1 vccd1 _13954_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12905_ _13100_/A _12905_/B vssd1 vssd1 vccd1 vccd1 _17922_/D sky130_fd_sc_hd__and2_1
X_16673_ _19246_/Q _16673_/B vssd1 vssd1 vccd1 vccd1 _16675_/B sky130_fd_sc_hd__nor2_1
XFILLER_262_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19461_ _19534_/CLK _19461_/D vssd1 vssd1 vccd1 vccd1 _19461_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_46_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13885_ _19325_/Q _13952_/A2 _13952_/B1 _13878_/X _13884_/X vssd1 vssd1 vccd1 vccd1
+ _13885_/Y sky130_fd_sc_hd__a2111oi_2
XFILLER_185_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18412_ _19591_/CLK _18412_/D vssd1 vssd1 vccd1 vccd1 _18412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15624_ _15789_/A1 _15619_/Y _15620_/X _15789_/B1 vssd1 vssd1 vccd1 vccd1 _15625_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ _12837_/A _12837_/B vssd1 vssd1 vccd1 vccd1 _12836_/Y sky130_fd_sc_hd__nor2_8
XFILLER_50_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _19526_/CLK _19392_/D vssd1 vssd1 vccd1 vccd1 _19392_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15555_ _15531_/A _15531_/B _15532_/A vssd1 vssd1 vccd1 vccd1 _15555_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18343_ _19621_/CLK _18343_/D vssd1 vssd1 vccd1 vccd1 _18343_/Q sky130_fd_sc_hd__dfxtp_1
X_12767_ _17824_/Q _13942_/A2 _13942_/B1 _17856_/Q vssd1 vssd1 vccd1 vccd1 _12767_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _16608_/A0 _18356_/Q _14517_/S vssd1 vssd1 vccd1 vccd1 _18356_/D sky130_fd_sc_hd__mux2_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18274_ _19231_/CLK _18274_/D vssd1 vssd1 vccd1 vccd1 _18274_/Q sky130_fd_sc_hd__dfxtp_1
X_11718_ _11919_/B _15835_/A _11968_/B2 vssd1 vssd1 vccd1 vccd1 _11718_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15486_ _15486_/A _15508_/B vssd1 vssd1 vccd1 vccd1 _15557_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12698_ _12697_/X _12696_/X _12818_/S vssd1 vssd1 vccd1 vccd1 _12698_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14437_ _18576_/Q _14451_/B vssd1 vssd1 vccd1 vccd1 _18289_/D sky130_fd_sc_hd__and2_1
X_17225_ _17223_/Y _17224_/X _17141_/A vssd1 vssd1 vccd1 vccd1 _19425_/D sky130_fd_sc_hd__a21oi_1
Xinput11 core_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_2
X_11649_ _11651_/B _11650_/B vssd1 vssd1 vccd1 vccd1 _11649_/Y sky130_fd_sc_hd__nor2_1
Xinput22 core_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
Xinput33 core_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17156_ _17255_/A _17156_/B vssd1 vssd1 vccd1 vccd1 _19403_/D sky130_fd_sc_hd__nor2_1
XFILLER_7_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 dout0[10] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_2
X_14368_ _18220_/Q _16542_/A0 _14377_/S vssd1 vssd1 vccd1 vccd1 _18220_/D sky130_fd_sc_hd__mux2_1
Xinput55 dout0[20] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_2
Xinput66 dout0[30] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput77 dout0[40] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_2
X_16107_ _18756_/Q _16137_/B vssd1 vssd1 vccd1 vccd1 _16107_/Y sky130_fd_sc_hd__nand2_1
Xinput88 dout0[50] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_2
X_13319_ _12442_/D _13315_/X _13318_/X vssd1 vssd1 vccd1 vccd1 _13319_/X sky130_fd_sc_hd__o21a_1
XFILLER_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput99 dout0[60] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_2
X_17087_ _19377_/Q _17107_/B vssd1 vssd1 vccd1 vccd1 _17087_/X sky130_fd_sc_hd__or2_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14299_ _16617_/A0 _18158_/Q _14305_/S vssd1 vssd1 vccd1 vccd1 _18158_/D sky130_fd_sc_hd__mux2_1
X_16038_ _16038_/A _16046_/A vssd1 vssd1 vccd1 vccd1 _18732_/D sky130_fd_sc_hd__and2_1
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_177_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18593_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08860_ input9/X vssd1 vssd1 vccd1 vccd1 _14528_/A sky130_fd_sc_hd__inv_2
XFILLER_111_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_106_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18761_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17989_ _18902_/CLK _17989_/D vssd1 vssd1 vccd1 vccd1 _17989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1890 _16128_/B1 vssd1 vssd1 vccd1 vccd1 _12187_/A sky130_fd_sc_hd__buf_2
XFILLER_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09412_ _10294_/A1 _19202_/Q _19170_/Q _09428_/B2 vssd1 vssd1 vccd1 vccd1 _09412_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_253_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09343_ _09341_/X _09342_/X _10169_/S vssd1 vssd1 vccd1 vccd1 _09343_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09274_ _09274_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _09274_/X sky130_fd_sc_hd__and2_1
XFILLER_178_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08989_ _11691_/B1 _12432_/A2 _08988_/X _11692_/A1 _18400_/Q vssd1 vssd1 vccd1 vccd1
+ _08999_/A sky130_fd_sc_hd__o32a_1
XFILLER_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10951_ _18255_/Q _18830_/Q _18458_/Q _18359_/Q _11340_/B2 _11357_/S1 vssd1 vssd1
+ vccd1 vccd1 _10952_/B sky130_fd_sc_hd__mux4_1
XFILLER_272_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13670_ _12733_/S _13194_/X _13669_/X vssd1 vssd1 vccd1 vccd1 _13670_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10882_ _11112_/A _10882_/B vssd1 vssd1 vccd1 vccd1 _10887_/A sky130_fd_sc_hd__and2_1
XFILLER_231_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12621_ _13225_/B _13225_/C _13225_/A vssd1 vssd1 vccd1 vccd1 _13226_/A sky130_fd_sc_hd__o21ai_2
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15340_ _15340_/A _15340_/B vssd1 vssd1 vccd1 vccd1 _15340_/Y sky130_fd_sc_hd__nor2_2
XFILLER_106_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12552_ _12552_/A _12552_/B vssd1 vssd1 vccd1 vccd1 _12552_/X sky130_fd_sc_hd__or2_2
XFILLER_240_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11503_ _18638_/Q _18060_/Q _19079_/Q _18983_/Q _11503_/S0 _11503_/S1 vssd1 vssd1
+ vccd1 vccd1 _11504_/B sky130_fd_sc_hd__mux4_1
XPHY_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15271_ _18570_/Q _15271_/B vssd1 vssd1 vccd1 vccd1 _15272_/B sky130_fd_sc_hd__nor2_1
X_12483_ _12483_/A _12483_/B vssd1 vssd1 vccd1 vccd1 _12483_/Y sky130_fd_sc_hd__nor2_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17010_ _17585_/A _17044_/A2 _17009_/X _17559_/A vssd1 vssd1 vccd1 vccd1 _19341_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14222_ _18109_/Q _14260_/B vssd1 vssd1 vccd1 vccd1 _14222_/X sky130_fd_sc_hd__or2_1
X_11434_ _11512_/A1 _19631_/Q _18920_/Q _11513_/B2 vssd1 vssd1 vccd1 vccd1 _11434_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14153_ _14153_/A _14153_/B _14153_/C _14153_/D vssd1 vssd1 vccd1 vccd1 _14158_/A
+ sky130_fd_sc_hd__and4_2
X_11365_ _11133_/B2 _11364_/X _11299_/X _11365_/B2 vssd1 vssd1 vccd1 vccd1 _15404_/A
+ sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_leaf_4_wb_clk_i _19652_/A vssd1 vssd1 vccd1 vccd1 _19600_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13104_ _19239_/Q _13425_/A2 _13425_/B1 _19271_/Q vssd1 vssd1 vccd1 vccd1 _13104_/X
+ sky130_fd_sc_hd__a22o_1
X_10316_ _19062_/Q _19030_/Q _10687_/S vssd1 vssd1 vccd1 vccd1 _10316_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14084_ _17667_/A0 _18024_/Q _14106_/S vssd1 vssd1 vccd1 vccd1 _18024_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18961_ _19602_/CLK _18961_/D vssd1 vssd1 vccd1 vccd1 _18961_/Q sky130_fd_sc_hd__dfxtp_1
X_11296_ _11219_/A _10086_/A _10679_/B _09039_/B vssd1 vssd1 vccd1 vccd1 _11296_/Y
+ sky130_fd_sc_hd__o22ai_1
X_17912_ _19595_/CLK _17912_/D vssd1 vssd1 vccd1 vccd1 _17912_/Q sky130_fd_sc_hd__dfxtp_4
X_13035_ _13349_/B _14142_/B vssd1 vssd1 vccd1 vccd1 _13035_/Y sky130_fd_sc_hd__nor2_1
X_10247_ _10243_/A _10246_/Y _10243_/Y _09264_/S vssd1 vssd1 vccd1 vccd1 _10247_/X
+ sky130_fd_sc_hd__a211o_1
X_18892_ _19635_/CLK _18892_/D vssd1 vssd1 vccd1 vccd1 _18892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1120 _13289_/A vssd1 vssd1 vccd1 vccd1 _13931_/A sky130_fd_sc_hd__buf_4
XFILLER_26_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1131 _12322_/Y vssd1 vssd1 vccd1 vccd1 _15416_/A sky130_fd_sc_hd__buf_6
X_17843_ _19470_/CLK _17843_/D vssd1 vssd1 vccd1 vccd1 _17843_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1142 _09859_/A vssd1 vssd1 vccd1 vccd1 _11333_/A1 sky130_fd_sc_hd__buf_8
X_10178_ _10176_/X _10177_/X _10253_/A vssd1 vssd1 vccd1 vccd1 _10178_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1153 _09079_/Y vssd1 vssd1 vccd1 vccd1 _13622_/A sky130_fd_sc_hd__buf_8
XFILLER_120_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1164 _15852_/X vssd1 vssd1 vccd1 vccd1 _15905_/C sky130_fd_sc_hd__buf_2
XFILLER_266_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1175 _14200_/S vssd1 vssd1 vccd1 vccd1 _14186_/S sky130_fd_sc_hd__buf_6
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1186 _10083_/X vssd1 vssd1 vccd1 vccd1 _11143_/A1 sky130_fd_sc_hd__buf_4
XFILLER_266_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1197 _15835_/X vssd1 vssd1 vccd1 vccd1 _16877_/B1 sky130_fd_sc_hd__buf_6
X_17774_ _19602_/CLK _17774_/D vssd1 vssd1 vccd1 vccd1 _17774_/Q sky130_fd_sc_hd__dfxtp_1
X_14986_ _14996_/A1 _14985_/X _15006_/B1 vssd1 vssd1 vccd1 vccd1 _14986_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_93_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19513_ _19546_/CLK _19513_/D vssd1 vssd1 vccd1 vccd1 _19513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16725_ _19261_/Q _16728_/C _12203_/A vssd1 vssd1 vccd1 vccd1 _16725_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13937_ _13937_/A _13937_/B vssd1 vssd1 vccd1 vccd1 _13937_/Y sky130_fd_sc_hd__nand2_1
XFILLER_208_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19444_ _19444_/CLK _19444_/D vssd1 vssd1 vccd1 vccd1 _19444_/Q sky130_fd_sc_hd__dfxtp_1
X_16656_ _19240_/Q _16658_/C _16655_/Y vssd1 vssd1 vccd1 vccd1 _19240_/D sky130_fd_sc_hd__o21a_1
X_13868_ _18129_/Q _13900_/C vssd1 vssd1 vccd1 vccd1 _13868_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_250_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12819_ _12728_/X _12734_/B _12821_/A vssd1 vssd1 vccd1 vccd1 _12933_/B sky130_fd_sc_hd__mux2_1
X_15607_ _19446_/Q _15793_/A2 _17202_/A _15606_/X vssd1 vssd1 vccd1 vccd1 _15607_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19375_ _19531_/CLK _19375_/D vssd1 vssd1 vccd1 vccd1 _19375_/Q sky130_fd_sc_hd__dfxtp_1
X_16587_ _17720_/A0 _19191_/Q _16589_/S vssd1 vssd1 vccd1 vccd1 _19191_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13799_ _12712_/S _13043_/Y _13048_/X _13863_/B2 _13798_/X vssd1 vssd1 vccd1 vccd1
+ _13799_/X sky130_fd_sc_hd__o221a_1
XFILLER_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18326_ _19573_/CLK _18326_/D vssd1 vssd1 vccd1 vccd1 _18326_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _15751_/A _15538_/B _15538_/C vssd1 vssd1 vccd1 vccd1 _15538_/X sky130_fd_sc_hd__or3_1
XFILLER_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18257_ _19639_/CLK _18257_/D vssd1 vssd1 vccd1 vccd1 _18257_/Q sky130_fd_sc_hd__dfxtp_1
X_15469_ _15369_/A _15464_/X _15468_/X _17540_/B1 vssd1 vssd1 vccd1 vccd1 _15469_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17208_ _17208_/A _17208_/B vssd1 vssd1 vccd1 vccd1 _17208_/Y sky130_fd_sc_hd__nand2_2
XFILLER_144_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18188_ _19641_/CLK _18188_/D vssd1 vssd1 vccd1 vccd1 _18188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _17157_/A _17571_/A vssd1 vssd1 vccd1 vccd1 _17423_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ _19619_/Q _18908_/Q _10281_/S vssd1 vssd1 vccd1 vccd1 _09961_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08912_ _17796_/Q _17794_/Q vssd1 vssd1 vccd1 vccd1 _08912_/Y sky130_fd_sc_hd__nor2_1
XFILLER_258_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _11131_/A _09886_/X _09889_/X _09891_/X _11279_/B1 vssd1 vssd1 vccd1 vccd1
+ _09892_/X sky130_fd_sc_hd__a311o_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08843_ _08843_/A vssd1 vssd1 vccd1 vccd1 _08843_/Y sky130_fd_sc_hd__inv_8
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_509 _10431_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18884_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_214_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09326_ _09326_/A _09326_/B vssd1 vssd1 vccd1 vccd1 _11141_/B sky130_fd_sc_hd__nor2_1
XFILLER_178_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09257_ _09255_/X _09256_/X _10409_/A vssd1 vssd1 vccd1 vccd1 _09257_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09188_ _11459_/B1 _09173_/X _09186_/X _09187_/X vssd1 vssd1 vccd1 vccd1 _09188_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ _11157_/A1 _19147_/Q _11160_/S _19115_/Q _09534_/S vssd1 vssd1 vccd1 vccd1
+ _11150_/X sky130_fd_sc_hd__o221a_1
XFILLER_1_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10101_ _18905_/Q _10101_/B vssd1 vssd1 vccd1 vccd1 _10101_/X sky130_fd_sc_hd__or2_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11081_ _10633_/A _11079_/X _11080_/X _11563_/B1 vssd1 vssd1 vccd1 vccd1 _11081_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput201 localMemory_wb_adr_i[1] vssd1 vssd1 vccd1 vccd1 input201/X sky130_fd_sc_hd__clkbuf_2
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput212 localMemory_wb_adr_i[8] vssd1 vssd1 vccd1 vccd1 input212/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10032_ _18594_/Q _18165_/Q _10500_/S vssd1 vssd1 vccd1 vccd1 _10032_/X sky130_fd_sc_hd__mux2_1
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput223 localMemory_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input223/X sky130_fd_sc_hd__clkbuf_16
XFILLER_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput234 localMemory_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 input234/X sky130_fd_sc_hd__clkbuf_16
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 localMemory_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input245/X sky130_fd_sc_hd__buf_8
Xinput256 manufacturerID[2] vssd1 vssd1 vccd1 vccd1 _15863_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput267 partID[12] vssd1 vssd1 vccd1 vccd1 input267/X sky130_fd_sc_hd__clkbuf_2
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _15003_/A1 _13436_/Y _15003_/B1 _18641_/Q _15003_/C1 vssd1 vssd1 vccd1 vccd1
+ _14840_/X sky130_fd_sc_hd__a221o_1
Xinput278 partID[8] vssd1 vssd1 vccd1 vccd1 _15914_/A sky130_fd_sc_hd__buf_2
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ _19228_/Q _15014_/B _14934_/C _14934_/D vssd1 vssd1 vccd1 vccd1 _14771_/X
+ sky130_fd_sc_hd__and4_4
X_11983_ _11980_/X _18725_/Q _15954_/B vssd1 vssd1 vccd1 vccd1 _11983_/X sky130_fd_sc_hd__mux2_1
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13722_ _19320_/Q _13754_/A2 _13722_/B1 _13715_/X _13721_/X vssd1 vssd1 vccd1 vccd1
+ _13722_/Y sky130_fd_sc_hd__a2111oi_2
X_16510_ _16543_/A0 _19116_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _19116_/D sky130_fd_sc_hd__mux2_1
X_10934_ _11584_/C1 _10931_/X _10932_/X _10933_/X vssd1 vssd1 vccd1 vccd1 _10934_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_216_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17490_ _13611_/B _17520_/A2 _17532_/A2 _17810_/Q _17538_/A vssd1 vssd1 vccd1 vccd1
+ _17490_/X sky130_fd_sc_hd__a221o_1
XFILLER_232_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16441_ _19049_/Q _17706_/A0 _16453_/S vssd1 vssd1 vccd1 vccd1 _19049_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ _19512_/Q _13947_/A2 _13781_/B1 _13652_/X vssd1 vssd1 vccd1 vccd1 _13653_/X
+ sky130_fd_sc_hd__o211a_1
X_10865_ _11584_/A1 _18153_/Q _18799_/Q _10864_/S vssd1 vssd1 vccd1 vccd1 _10865_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12604_ _12842_/A _12842_/B vssd1 vssd1 vccd1 vccd1 _12604_/Y sky130_fd_sc_hd__nand2_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19160_ _19613_/CLK _19160_/D vssd1 vssd1 vccd1 vccd1 _19160_/Q sky130_fd_sc_hd__dfxtp_1
X_16372_ _17704_/A0 _18983_/Q _16390_/S vssd1 vssd1 vccd1 vccd1 _18983_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _19252_/Q _13625_/A2 _13625_/B1 _19284_/Q vssd1 vssd1 vccd1 vccd1 _13584_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_158_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10796_ _18553_/Q _18428_/Q _11604_/S vssd1 vssd1 vccd1 vccd1 _10796_/X sky130_fd_sc_hd__mux2_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _18741_/CLK _18111_/D vssd1 vssd1 vccd1 vccd1 _18111_/Q sky130_fd_sc_hd__dfxtp_4
X_15323_ _19465_/Q _19399_/Q _15322_/X vssd1 vssd1 vccd1 vccd1 _15324_/B sky130_fd_sc_hd__o21ai_2
X_12535_ _12577_/A _13165_/B vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__or2_4
XFILLER_169_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19091_ _19155_/CLK _19091_/D vssd1 vssd1 vccd1 vccd1 _19091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18042_ _19612_/CLK _18042_/D vssd1 vssd1 vccd1 vccd1 _18042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15254_ _15254_/A _15254_/B vssd1 vssd1 vccd1 vccd1 _15254_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_184_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12466_ _12466_/A0 _14672_/C _12482_/S vssd1 vssd1 vccd1 vccd1 _12513_/B sky130_fd_sc_hd__mux2_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14205_ _14205_/A _14205_/B vssd1 vssd1 vccd1 vccd1 _18100_/D sky130_fd_sc_hd__and2_1
XFILLER_126_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11417_ _11428_/A _11416_/X _11417_/B1 vssd1 vssd1 vccd1 vccd1 _11417_/X sky130_fd_sc_hd__a21o_1
XFILLER_137_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15185_ _15167_/A _15166_/B _15166_/A vssd1 vssd1 vccd1 vccd1 _15189_/A sky130_fd_sc_hd__o21ba_1
X_12397_ _12427_/A _12397_/B vssd1 vssd1 vccd1 vccd1 _12397_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14136_ _16553_/A0 _18075_/Q _14139_/S vssd1 vssd1 vccd1 vccd1 _18075_/D sky130_fd_sc_hd__mux2_1
XFILLER_235_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11348_ _11358_/A _11347_/X _11608_/C1 vssd1 vssd1 vccd1 vccd1 _11348_/X sky130_fd_sc_hd__a21o_1
XFILLER_113_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18944_ _19211_/CLK _18944_/D vssd1 vssd1 vccd1 vccd1 _18944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14067_ _16551_/A0 _18009_/Q _14073_/S vssd1 vssd1 vccd1 vccd1 _18009_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11279_ _10745_/S _11278_/X _11279_/B1 vssd1 vssd1 vccd1 vccd1 _11280_/B sky130_fd_sc_hd__a21o_1
XFILLER_279_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13018_ _19333_/Q _13246_/A2 _13246_/B1 _19461_/Q _12570_/C vssd1 vssd1 vccd1 vccd1
+ _13018_/X sky130_fd_sc_hd__a221o_1
X_18875_ _18875_/CLK _18875_/D vssd1 vssd1 vccd1 vccd1 _18875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_255_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17826_ _18713_/CLK _17826_/D vssd1 vssd1 vccd1 vccd1 _17826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17757_ _18657_/Q vssd1 vssd1 vccd1 vccd1 _18657_/D sky130_fd_sc_hd__clkbuf_2
X_14969_ _14979_/A1 _18272_/Q _14968_/Y _11712_/A vssd1 vssd1 vccd1 vccd1 _14969_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16708_ _19255_/Q _19254_/Q _19253_/Q _16708_/D vssd1 vssd1 vccd1 vccd1 _16717_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_63_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17688_ _17688_/A0 _19615_/Q _17689_/S vssd1 vssd1 vccd1 vccd1 _19615_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19427_ _19507_/CLK _19427_/D vssd1 vssd1 vccd1 vccd1 _19427_/Q sky130_fd_sc_hd__dfxtp_1
X_16639_ _16752_/A _16639_/B _16643_/C vssd1 vssd1 vccd1 vccd1 _19235_/D sky130_fd_sc_hd__nor3_1
XFILLER_250_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19358_ _19458_/CLK _19358_/D vssd1 vssd1 vccd1 vccd1 _19358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09111_ _18854_/Q _11167_/B _09845_/S _09110_/X vssd1 vssd1 vccd1 vccd1 _09111_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_149_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18309_ _19620_/CLK _18309_/D vssd1 vssd1 vccd1 vccd1 _18309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19289_ _19291_/CLK _19289_/D vssd1 vssd1 vccd1 vccd1 _19289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09042_ _09042_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _09042_/Y sky130_fd_sc_hd__nand2_2
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_192_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19642_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_121_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19310_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout902 _16204_/A0 vssd1 vssd1 vccd1 vccd1 _16535_/A0 sky130_fd_sc_hd__clkbuf_4
X_09944_ _15120_/A _11785_/B _09943_/Y _09697_/B vssd1 vssd1 vccd1 vccd1 _09944_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout913 _16359_/X vssd1 vssd1 vccd1 vccd1 _16385_/S sky130_fd_sc_hd__buf_12
Xfanout924 _16212_/S vssd1 vssd1 vccd1 vccd1 _16226_/S sky130_fd_sc_hd__buf_12
Xfanout935 _14679_/X vssd1 vssd1 vccd1 vccd1 _14983_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout946 _14670_/Y vssd1 vssd1 vccd1 vccd1 _14913_/B1 sky130_fd_sc_hd__buf_2
XFILLER_258_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout957 _14521_/S vssd1 vssd1 vccd1 vccd1 _14516_/S sky130_fd_sc_hd__buf_12
X_09875_ _10036_/S _09873_/X _09874_/X _10589_/S vssd1 vssd1 vccd1 vccd1 _09875_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout968 _14075_/Y vssd1 vssd1 vccd1 vccd1 _14104_/S sky130_fd_sc_hd__buf_12
XFILLER_258_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout979 _12463_/X vssd1 vssd1 vccd1 vccd1 _13115_/B2 sky130_fd_sc_hd__buf_4
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _18740_/Q vssd1 vssd1 vccd1 vccd1 _11981_/B sky130_fd_sc_hd__inv_2
XFILLER_245_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_306 _18113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_317 _18128_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_328 _11959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_339 _11482_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10650_ _19090_/Q _18994_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _10650_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09309_ _09967_/S _09302_/X _09301_/X _11507_/S vssd1 vssd1 vccd1 vccd1 _09309_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10581_ _18260_/Q _18835_/Q _10582_/S vssd1 vssd1 vccd1 vccd1 _10581_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12320_ _12320_/A _12320_/B _12320_/C _11482_/A2 vssd1 vssd1 vccd1 vccd1 _12321_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_155_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ _16808_/A _12251_/B vssd1 vssd1 vccd1 vccd1 _12251_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11202_ _18548_/Q _18423_/Q _18032_/Q _18000_/Q _10726_/S _11274_/S1 vssd1 vssd1
+ vccd1 vccd1 _11202_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _17857_/Q _12184_/C _12181_/Y vssd1 vssd1 vccd1 vccd1 _17857_/D sky130_fd_sc_hd__o21a_1
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11133_ _11365_/B2 _11067_/X _11132_/X _11133_/B2 vssd1 vssd1 vccd1 vccd1 _15478_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16990_ _19331_/Q _17043_/B _16989_/Y _17378_/A vssd1 vssd1 vccd1 vccd1 _19331_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15941_ input6/X _12770_/A _15941_/S vssd1 vssd1 vccd1 vccd1 _15941_/X sky130_fd_sc_hd__mux2_1
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11064_ _09574_/A _09239_/X _11064_/B1 vssd1 vssd1 vccd1 vccd1 _11066_/A sky130_fd_sc_hd__a21oi_1
XFILLER_150_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10015_ _10013_/X _10014_/X _11568_/A vssd1 vssd1 vccd1 vccd1 _10015_/X sky130_fd_sc_hd__mux2_1
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _18660_/CLK _18660_/D vssd1 vssd1 vccd1 vccd1 _18660_/Q sky130_fd_sc_hd__dfxtp_1
X_15872_ _15872_/A _15881_/B _15908_/C vssd1 vssd1 vccd1 vccd1 _15872_/X sky130_fd_sc_hd__and3_1
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17611_ _15093_/C _17592_/X _17623_/B1 vssd1 vssd1 vccd1 vccd1 _17611_/X sky130_fd_sc_hd__a21o_1
XFILLER_264_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ _15006_/A1 _14822_/X _14875_/B1 vssd1 vssd1 vccd1 vccd1 _14823_/Y sky130_fd_sc_hd__o21ai_2
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _19453_/CLK _18591_/D vssd1 vssd1 vccd1 vccd1 _18591_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_224_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _19519_/Q _17493_/B _17541_/X vssd1 vssd1 vccd1 vccd1 _19519_/D sky130_fd_sc_hd__o21ba_1
X_14754_ _14865_/A1 _14753_/X _14865_/B1 vssd1 vssd1 vccd1 vccd1 _14754_/Y sky130_fd_sc_hd__o21ai_2
X_11966_ _18512_/Q _11720_/X _11916_/X _11968_/B2 vssd1 vssd1 vccd1 vccd1 _11966_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_217_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ _18123_/Q _13704_/C _18124_/Q vssd1 vssd1 vccd1 vccd1 _13706_/B sky130_fd_sc_hd__a21oi_1
X_10917_ _11562_/S _10916_/X _10915_/X _11084_/S vssd1 vssd1 vccd1 vccd1 _10917_/X
+ sky130_fd_sc_hd__a211o_1
X_14685_ _19227_/Q _14934_/C vssd1 vssd1 vccd1 vccd1 _14685_/X sky130_fd_sc_hd__and2_1
X_17473_ _17473_/A _17493_/B vssd1 vssd1 vccd1 vccd1 _17473_/Y sky130_fd_sc_hd__nand2_1
X_11897_ _11823_/A _11832_/B _11875_/A _11896_/X vssd1 vssd1 vccd1 vccd1 _11897_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_232_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19212_ _19621_/CLK _19212_/D vssd1 vssd1 vccd1 vccd1 _19212_/Q sky130_fd_sc_hd__dfxtp_1
X_16424_ _16490_/A0 _19033_/Q _16424_/S vssd1 vssd1 vccd1 vccd1 _19033_/D sky130_fd_sc_hd__mux2_1
XFILLER_220_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13636_ _14016_/B vssd1 vssd1 vccd1 vccd1 _13636_/Y sky130_fd_sc_hd__inv_2
X_10848_ _11311_/C1 _10847_/X _10846_/X _11577_/S vssd1 vssd1 vccd1 vccd1 _10848_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19143_ _19157_/CLK _19143_/D vssd1 vssd1 vccd1 vccd1 _19143_/Q sky130_fd_sc_hd__dfxtp_1
X_16355_ _18967_/Q _16488_/A0 _16355_/S vssd1 vssd1 vccd1 vccd1 _18967_/D sky130_fd_sc_hd__mux2_1
X_13567_ _12593_/A _13533_/B _12594_/X vssd1 vssd1 vccd1 vccd1 _13568_/B sky130_fd_sc_hd__o21ai_2
XFILLER_201_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10779_ _10777_/X _10778_/X _10784_/S vssd1 vssd1 vccd1 vccd1 _10779_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12518_ _12554_/A _12554_/B _12512_/B vssd1 vssd1 vccd1 vccd1 _12577_/B sky130_fd_sc_hd__or3b_4
XFILLER_9_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15306_ _12442_/A _15113_/Y _15305_/X vssd1 vssd1 vccd1 vccd1 _15306_/Y sky130_fd_sc_hd__a21oi_1
X_19074_ _19138_/CLK _19074_/D vssd1 vssd1 vccd1 vccd1 _19074_/Q sky130_fd_sc_hd__dfxtp_1
X_16286_ _17717_/A0 _18900_/Q _16292_/S vssd1 vssd1 vccd1 vccd1 _18900_/D sky130_fd_sc_hd__mux2_1
X_13498_ _19507_/Q _13781_/A2 _13781_/B1 _13497_/X vssd1 vssd1 vccd1 vccd1 _13498_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18025_ _19595_/CLK _18025_/D vssd1 vssd1 vccd1 vccd1 _18025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12449_ _13421_/A _13462_/A _15083_/A _12461_/A vssd1 vssd1 vccd1 vccd1 _12449_/X
+ sky130_fd_sc_hd__o31a_2
X_15237_ _18568_/Q _15447_/B _15235_/X _15236_/Y _14430_/B vssd1 vssd1 vccd1 vccd1
+ _18568_/D sky130_fd_sc_hd__o221a_1
XFILLER_160_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15168_ _19459_/Q _15167_/Y _15400_/S vssd1 vssd1 vccd1 vccd1 _15168_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14119_ _16470_/A0 _18058_/Q _14139_/S vssd1 vssd1 vccd1 vccd1 _18058_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15099_ _19389_/Q _15092_/B input175/X _15092_/X vssd1 vssd1 vccd1 vccd1 _15099_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_262_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18927_ _19638_/CLK _18927_/D vssd1 vssd1 vccd1 vccd1 _18927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_268_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09660_ _10085_/A _09660_/B _09660_/C vssd1 vssd1 vccd1 vccd1 _09660_/X sky130_fd_sc_hd__or3_2
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18858_ _19601_/CLK _18858_/D vssd1 vssd1 vccd1 vccd1 _18858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17809_ _17814_/CLK _17809_/D vssd1 vssd1 vccd1 vccd1 _17809_/Q sky130_fd_sc_hd__dfxtp_4
X_09591_ _09579_/X _09590_/X _10746_/S vssd1 vssd1 vccd1 vccd1 _09591_/X sky130_fd_sc_hd__mux2_1
XFILLER_282_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18789_ _19203_/CLK _18789_/D vssd1 vssd1 vccd1 vccd1 _18789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_283_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XExperiarCore_1911 vssd1 vssd1 vccd1 vccd1 ExperiarCore_1911/HI localMemory_wb_error_o
+ sky130_fd_sc_hd__conb_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ _09025_/A _09025_/B vssd1 vssd1 vccd1 vccd1 _09048_/A sky130_fd_sc_hd__nand2_4
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout710 _13115_/C1 vssd1 vssd1 vccd1 vccd1 _13854_/B1 sky130_fd_sc_hd__buf_4
Xfanout1708 _09750_/S vssd1 vssd1 vccd1 vccd1 _11578_/S sky130_fd_sc_hd__buf_8
XFILLER_278_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout721 _12497_/Y vssd1 vssd1 vccd1 vccd1 _13844_/B1 sky130_fd_sc_hd__buf_4
XFILLER_172_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1719 _19231_/Q vssd1 vssd1 vccd1 vccd1 _12461_/A sky130_fd_sc_hd__buf_12
XFILLER_131_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout732 _16539_/A0 vssd1 vssd1 vccd1 vccd1 _17705_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09927_ _09845_/S _09925_/X _09926_/X vssd1 vssd1 vccd1 vccd1 _09927_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout743 _11223_/X vssd1 vssd1 vccd1 vccd1 _17641_/A0 sky130_fd_sc_hd__clkbuf_8
Xfanout754 _12609_/A vssd1 vssd1 vccd1 vccd1 _13390_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout765 _17723_/S vssd1 vssd1 vccd1 vccd1 _17718_/S sky130_fd_sc_hd__buf_12
Xfanout776 _17625_/Y vssd1 vssd1 vccd1 vccd1 _17654_/S sky130_fd_sc_hd__buf_12
Xfanout787 _16554_/S vssd1 vssd1 vccd1 vccd1 _16556_/S sky130_fd_sc_hd__buf_12
X_09858_ _09849_/X _09857_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09859_/C sky130_fd_sc_hd__o21ai_2
XFILLER_246_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout798 _16325_/S vssd1 vssd1 vccd1 vccd1 _16323_/S sky130_fd_sc_hd__buf_12
XFILLER_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _10589_/S _09789_/B vssd1 vssd1 vccd1 vccd1 _09789_/Y sky130_fd_sc_hd__nor2_1
XFILLER_283_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11820_/A _11820_/B vssd1 vssd1 vccd1 vccd1 _11820_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_103 _11819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _11807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _11865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _11831_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _11868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11751_/A vssd1 vssd1 vccd1 vccd1 _11751_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_158 _11909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_169 _13141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _10315_/S _10701_/X _11237_/B1 vssd1 vssd1 vccd1 vccd1 _10702_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _18322_/Q _17674_/A0 _14477_/S vssd1 vssd1 vccd1 vccd1 _18322_/D sky130_fd_sc_hd__mux2_1
X_11682_ _13330_/B vssd1 vssd1 vccd1 vccd1 _11683_/B sky130_fd_sc_hd__inv_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13421_ _13421_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _13421_/Y sky130_fd_sc_hd__nand2_1
X_10633_ _10633_/A _10633_/B vssd1 vssd1 vccd1 vccd1 _10633_/X sky130_fd_sc_hd__or2_1
X_16140_ _16140_/A1 _16139_/Y _16142_/B1 vssd1 vssd1 vccd1 vccd1 _18772_/D sky130_fd_sc_hd__a21oi_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13352_ _13312_/A _14145_/A _13909_/B1 vssd1 vssd1 vccd1 vccd1 _13352_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10564_ _11103_/A _10564_/B vssd1 vssd1 vccd1 vccd1 _10564_/Y sky130_fd_sc_hd__nor2_1
X_12303_ _18100_/Q _18099_/Q _18098_/Q vssd1 vssd1 vccd1 vccd1 _12303_/X sky130_fd_sc_hd__or3_4
XFILLER_6_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16071_ _16075_/A _16068_/X _16070_/Y _16053_/Y vssd1 vssd1 vccd1 vccd1 _16071_/Y
+ sky130_fd_sc_hd__a211oi_1
X_13283_ _19307_/Q _12583_/Y _13281_/X _13282_/X vssd1 vssd1 vccd1 vccd1 _13283_/X
+ sky130_fd_sc_hd__a211o_1
X_10495_ _18041_/Q _18009_/Q _10500_/S vssd1 vssd1 vccd1 vccd1 _10495_/X sky130_fd_sc_hd__mux2_1
X_15022_ _18511_/Q input211/X _15024_/S vssd1 vssd1 vccd1 vccd1 _18511_/D sky130_fd_sc_hd__mux2_1
X_12234_ _17877_/Q _12234_/B vssd1 vssd1 vccd1 vccd1 _12240_/C sky130_fd_sc_hd__and2_2
XFILLER_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12165_ _17851_/Q _12168_/C _16808_/A vssd1 vssd1 vccd1 vccd1 _12165_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_268_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11116_ _10040_/S _11115_/X _11623_/A1 vssd1 vssd1 vccd1 vccd1 _11117_/B sky130_fd_sc_hd__a21o_1
XFILLER_123_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12096_ _12107_/A _12096_/B _12100_/C vssd1 vssd1 vccd1 vccd1 _17825_/D sky130_fd_sc_hd__nor3_1
X_16973_ _17118_/B _16973_/B vssd1 vssd1 vccd1 vccd1 _17555_/B sky130_fd_sc_hd__or2_4
XFILLER_111_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18712_ _18713_/CLK _18712_/D vssd1 vssd1 vccd1 vccd1 _18712_/Q sky130_fd_sc_hd__dfxtp_1
X_15924_ _18683_/Q _15948_/A2 _15945_/C1 _15923_/X vssd1 vssd1 vccd1 vccd1 _15924_/X
+ sky130_fd_sc_hd__a211o_1
X_11047_ _11512_/A1 _19604_/Q _19572_/Q _11426_/B2 vssd1 vssd1 vccd1 vccd1 _11047_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 core_wb_ack_i vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18643_ _19586_/CLK _18643_/D vssd1 vssd1 vccd1 vccd1 _18643_/Q sky130_fd_sc_hd__dfxtp_4
X_15855_ _15854_/A _16002_/A2 _15908_/C _18735_/Q _15906_/B1 vssd1 vssd1 vccd1 vccd1
+ _15855_/X sky130_fd_sc_hd__a221o_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _14696_/A _18270_/Q _14805_/Y _14846_/B1 vssd1 vssd1 vccd1 vccd1 _14806_/X
+ sky130_fd_sc_hd__a31o_1
X_18574_ _19531_/CLK _18574_/D vssd1 vssd1 vccd1 vccd1 _18574_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ _14268_/A _15786_/A2 _15785_/X _15481_/B vssd1 vssd1 vccd1 vccd1 _15787_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_280_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _12992_/Y _12997_/Y _13315_/S vssd1 vssd1 vccd1 vccd1 _12998_/X sky130_fd_sc_hd__mux2_2
XFILLER_252_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ _17817_/Q _17532_/A2 _17531_/B _13810_/A vssd1 vssd1 vccd1 vccd1 _17525_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_91_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14737_ input87/X input72/X _14784_/S vssd1 vssd1 vccd1 vccd1 _14737_/X sky130_fd_sc_hd__mux2_8
X_11949_ _14667_/A1 _11899_/B _11899_/C _11949_/B1 input236/X vssd1 vssd1 vccd1 vccd1
+ _11949_/X sky130_fd_sc_hd__a32o_4
XFILLER_221_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17456_ _18575_/Q _17461_/A2 _17455_/X _17546_/A2 vssd1 vssd1 vccd1 vccd1 _17456_/X
+ sky130_fd_sc_hd__o211a_1
X_14668_ _14688_/A _14669_/B vssd1 vssd1 vccd1 vccd1 _14681_/B sky130_fd_sc_hd__nor2_1
XFILLER_220_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16407_ _11376_/B _19016_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _19016_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _13616_/A _12265_/B _13618_/X vssd1 vssd1 vccd1 vccd1 _13619_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_220_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17387_ _17386_/B _17428_/A _17382_/A _19488_/Q vssd1 vssd1 vccd1 vccd1 _17387_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_14599_ _14599_/A _16359_/A vssd1 vssd1 vccd1 vccd1 _14599_/X sky130_fd_sc_hd__or2_4
XFILLER_220_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19126_ _19126_/CLK _19126_/D vssd1 vssd1 vccd1 vccd1 _19126_/Q sky130_fd_sc_hd__dfxtp_1
X_16338_ _18950_/Q _17670_/A0 _16357_/S vssd1 vssd1 vccd1 vccd1 _18950_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19057_ _19623_/CLK _19057_/D vssd1 vssd1 vccd1 vccd1 _19057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16269_ _17700_/A0 _18883_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _18883_/D sky130_fd_sc_hd__mux2_1
XFILLER_195_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput302 _11918_/X vssd1 vssd1 vccd1 vccd1 addr1[8] sky130_fd_sc_hd__buf_4
X_18008_ _19638_/CLK _18008_/D vssd1 vssd1 vccd1 vccd1 _18008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput313 _11761_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[17] sky130_fd_sc_hd__buf_4
Xoutput324 _11771_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[27] sky130_fd_sc_hd__buf_4
Xoutput335 _11814_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[10] sky130_fd_sc_hd__buf_4
Xoutput346 _11857_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[20] sky130_fd_sc_hd__buf_4
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput357 _11904_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[30] sky130_fd_sc_hd__buf_4
XFILLER_259_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput368 _11778_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[2] sky130_fd_sc_hd__buf_4
XFILLER_273_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput379 _11932_/X vssd1 vssd1 vccd1 vccd1 din0[12] sky130_fd_sc_hd__buf_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09712_ _19622_/Q _18911_/Q _09720_/S vssd1 vssd1 vccd1 vccd1 _09712_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09643_ _09643_/A _11796_/B vssd1 vssd1 vccd1 vccd1 _09643_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _09574_/A _09574_/B _09574_/C vssd1 vssd1 vccd1 vccd1 _09574_/X sky130_fd_sc_hd__or3_2
XFILLER_270_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09008_ input122/X input157/X _09655_/S vssd1 vssd1 vccd1 vccd1 _09008_/X sky130_fd_sc_hd__mux2_8
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10280_ _10278_/X _10279_/X _10280_/S vssd1 vssd1 vccd1 vccd1 _10280_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1505 fanout1525/X vssd1 vssd1 vccd1 vccd1 _08968_/S0 sky130_fd_sc_hd__buf_4
Xfanout1516 fanout1524/X vssd1 vssd1 vccd1 vccd1 _09290_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_278_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1527 _10643_/S vssd1 vssd1 vccd1 vccd1 _11112_/A sky130_fd_sc_hd__buf_6
XFILLER_265_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1538 _09967_/S vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__buf_6
Xfanout540 _15126_/X vssd1 vssd1 vccd1 vccd1 _15633_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout551 _17202_/A vssd1 vssd1 vccd1 vccd1 _17214_/A sky130_fd_sc_hd__buf_8
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1549 _08899_/Y vssd1 vssd1 vccd1 vccd1 _10033_/S sky130_fd_sc_hd__buf_6
XFILLER_247_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout562 _15437_/B1 vssd1 vssd1 vccd1 vccd1 _15307_/B sky130_fd_sc_hd__buf_6
Xfanout573 _16142_/A1 vssd1 vssd1 vccd1 vccd1 _16140_/A1 sky130_fd_sc_hd__buf_4
X_13970_ _15452_/A _13968_/X _13969_/Y _13970_/B2 vssd1 vssd1 vccd1 vccd1 _13970_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_281_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout584 _12024_/Y vssd1 vssd1 vccd1 vccd1 _12052_/A2 sky130_fd_sc_hd__buf_4
XFILLER_281_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout595 _14268_/B vssd1 vssd1 vccd1 vccd1 _14252_/B sky130_fd_sc_hd__buf_4
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _13303_/B2 _12907_/X _12920_/X vssd1 vssd1 vccd1 vccd1 _13980_/B sky130_fd_sc_hd__a21oi_4
XFILLER_234_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15640_ _15787_/A _15640_/B vssd1 vssd1 vccd1 vccd1 _15640_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12852_ _19524_/Q _19492_/Q _13277_/S vssd1 vssd1 vccd1 vccd1 _12852_/X sky130_fd_sc_hd__mux2_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _11820_/A _11803_/B vssd1 vssd1 vccd1 vccd1 _11803_/Y sky130_fd_sc_hd__nor2_2
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _13115_/B2 _12767_/X _12782_/X vssd1 vssd1 vccd1 vccd1 _13976_/B sky130_fd_sc_hd__a21oi_4
X_15571_ _19476_/Q _15570_/X _15781_/S vssd1 vssd1 vccd1 vccd1 _15571_/X sky130_fd_sc_hd__mux2_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17310_ _19454_/Q _17310_/B vssd1 vssd1 vccd1 vccd1 _17310_/Y sky130_fd_sc_hd__nand2_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14522_ _14244_/B _14522_/A2 _11818_/B vssd1 vssd1 vccd1 vccd1 _14522_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11734_/A _11734_/B vssd1 vssd1 vccd1 vccd1 _12957_/A sky130_fd_sc_hd__nor2_8
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18290_ _19453_/CLK _18290_/D vssd1 vssd1 vccd1 vccd1 _18290_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _19431_/Q _17241_/B vssd1 vssd1 vccd1 vccd1 _17241_/Y sky130_fd_sc_hd__nand2_1
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14453_ _18593_/Q _17356_/A vssd1 vssd1 vccd1 vccd1 _18306_/D sky130_fd_sc_hd__and2_1
X_11665_ _18573_/Q _11663_/A _13258_/A _11664_/X vssd1 vssd1 vccd1 vccd1 _11704_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_168_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13404_ _17934_/Q _13742_/A2 _13403_/X _14181_/A vssd1 vssd1 vccd1 vccd1 _17934_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10616_ _18259_/Q _18834_/Q _10619_/S vssd1 vssd1 vccd1 vccd1 _10616_/X sky130_fd_sc_hd__mux2_1
X_14384_ _16459_/A _16459_/B _16194_/B _14074_/B vssd1 vssd1 vccd1 vccd1 _14384_/X
+ sky130_fd_sc_hd__or4b_4
X_17172_ _17211_/A _17172_/B vssd1 vssd1 vccd1 vccd1 _17478_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11596_ _11596_/A1 _18164_/Q _18810_/Q _10815_/B _08899_/A vssd1 vssd1 vccd1 vccd1
+ _11596_/X sky130_fd_sc_hd__a221o_1
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13335_ _19245_/Q _13495_/A2 _13495_/B1 _19277_/Q vssd1 vssd1 vccd1 vccd1 _13335_/X
+ sky130_fd_sc_hd__a22o_1
X_16123_ _18764_/Q _16139_/B vssd1 vssd1 vccd1 vccd1 _16123_/Y sky130_fd_sc_hd__nand2_1
X_10547_ _18157_/Q _11482_/A2 _10546_/X _11578_/S vssd1 vssd1 vccd1 vccd1 _10547_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_41_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16054_ _16054_/A _16069_/A vssd1 vssd1 vccd1 vccd1 _16055_/A sky130_fd_sc_hd__or2_2
X_13266_ _13315_/S _12992_/Y _13413_/B1 vssd1 vssd1 vccd1 vccd1 _13266_/X sky130_fd_sc_hd__a21o_2
XFILLER_142_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10478_ _10707_/A _10477_/X _11563_/B1 vssd1 vssd1 vccd1 vccd1 _10478_/X sky130_fd_sc_hd__o21a_1
X_12217_ _12219_/A _12217_/B _12218_/B vssd1 vssd1 vccd1 vccd1 _17870_/D sky130_fd_sc_hd__nor3_1
XFILLER_170_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15005_ _18132_/Q _14893_/S _14934_/X _15004_/X vssd1 vssd1 vccd1 vccd1 _15005_/X
+ sky130_fd_sc_hd__o211a_2
X_13197_ _13194_/S _13091_/X _13197_/B1 vssd1 vssd1 vccd1 vccd1 _13197_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12148_ _17844_/Q _12146_/B _12147_/Y vssd1 vssd1 vccd1 vccd1 _17844_/D sky130_fd_sc_hd__o21a_1
XFILLER_257_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16956_ _16960_/A _16956_/B vssd1 vssd1 vccd1 vccd1 _19323_/D sky130_fd_sc_hd__and2_1
X_12079_ _17817_/Q _12085_/B vssd1 vssd1 vccd1 vccd1 _12079_/X sky130_fd_sc_hd__or2_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15907_ _18678_/Q _15910_/A2 _15906_/X _15910_/C1 vssd1 vssd1 vccd1 vccd1 _18678_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16887_ _19306_/Q _17579_/A _16971_/S vssd1 vssd1 vccd1 vccd1 _16888_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18626_ _19197_/CLK _18626_/D vssd1 vssd1 vccd1 vccd1 _18626_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_266_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _18658_/Q _15843_/A _15837_/Y _17322_/A vssd1 vssd1 vccd1 vccd1 _18658_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18557_ _19092_/CLK _18557_/D vssd1 vssd1 vccd1 vccd1 _18557_/Q sky130_fd_sc_hd__dfxtp_1
X_15769_ _15728_/A _15728_/B _15749_/A _15768_/Y vssd1 vssd1 vccd1 vccd1 _15770_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17508_ _17508_/A _17517_/B vssd1 vssd1 vccd1 vccd1 _17508_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09290_ _19044_/Q _19012_/Q _09290_/S vssd1 vssd1 vccd1 vccd1 _09290_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18488_ _19286_/CLK _18488_/D vssd1 vssd1 vccd1 vccd1 _18488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_14 _14869_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ _19499_/Q _17547_/B _17437_/X _17438_/Y _17469_/C1 vssd1 vssd1 vccd1 vccd1
+ _19499_/D sky130_fd_sc_hd__o221a_1
XANTENNA_25 _15955_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_36 _09045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_47 _12612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_58 _11785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_69 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19109_ _19604_/CLK _19109_/D vssd1 vssd1 vccd1 vccd1 _19109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_99_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19079_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_28_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18201_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_161_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09626_ _11173_/S _09625_/X _09624_/X vssd1 vssd1 vccd1 vccd1 _09626_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09557_ _09611_/A _15808_/A1 _09556_/Y vssd1 vssd1 vccd1 vccd1 _11798_/B sky130_fd_sc_hd__o21ai_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09488_ _09027_/A _09034_/B _09487_/X _10084_/B _09483_/Y vssd1 vssd1 vccd1 vccd1
+ _09489_/C sky130_fd_sc_hd__a32o_1
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ _09987_/A _11449_/X _11447_/X vssd1 vssd1 vccd1 vccd1 _11450_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10401_ _11465_/A1 _19580_/Q _11462_/S _19612_/Q vssd1 vssd1 vccd1 vccd1 _10401_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11381_ _11465_/A1 _18217_/Q _11384_/B _18952_/Q _11464_/C1 vssd1 vssd1 vccd1 vccd1
+ _11381_/X sky130_fd_sc_hd__o221a_1
XFILLER_165_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _13438_/A _13101_/Y _13563_/B1 vssd1 vssd1 vccd1 vccd1 _13120_/X sky130_fd_sc_hd__a21o_1
X_10332_ _10338_/A1 _10327_/X _10331_/X vssd1 vssd1 vccd1 vccd1 _10332_/X sky130_fd_sc_hd__o21a_2
XFILLER_164_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _13051_/A _13051_/B _13051_/C vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__or3_1
X_10263_ _10263_/A1 _19159_/Q _09937_/S _19127_/Q vssd1 vssd1 vccd1 vccd1 _10263_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12002_ _17769_/Q _17703_/A0 _12021_/S vssd1 vssd1 vccd1 vccd1 _17769_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1302 _16961_/A2 vssd1 vssd1 vccd1 vccd1 _16969_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_267_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10194_ _10180_/A _10193_/Y _10180_/Y _10194_/C1 vssd1 vssd1 vccd1 vccd1 _10194_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1313 _11724_/Y vssd1 vssd1 vccd1 vccd1 _14349_/B sky130_fd_sc_hd__buf_6
XFILLER_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1324 _09098_/Y vssd1 vssd1 vccd1 vccd1 _11563_/B1 sky130_fd_sc_hd__clkbuf_16
X_16810_ _19292_/Q _16810_/B vssd1 vssd1 vccd1 vccd1 _16815_/C sky130_fd_sc_hd__and2_2
Xfanout1335 _11459_/A1 vssd1 vssd1 vccd1 vccd1 _10169_/S sky130_fd_sc_hd__buf_6
Xfanout1346 _10841_/C1 vssd1 vssd1 vccd1 vccd1 _09853_/S sky130_fd_sc_hd__buf_8
X_17790_ _19650_/CLK _17790_/D vssd1 vssd1 vccd1 vccd1 _17790_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1357 _10838_/B vssd1 vssd1 vccd1 vccd1 _11300_/B sky130_fd_sc_hd__buf_6
XFILLER_238_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1368 _10929_/S vssd1 vssd1 vccd1 vccd1 _10853_/S sky130_fd_sc_hd__buf_6
Xfanout1379 _11073_/B1 vssd1 vssd1 vccd1 vccd1 _11581_/S sky130_fd_sc_hd__buf_6
X_16741_ _19266_/Q _16743_/C _16740_/Y vssd1 vssd1 vccd1 vccd1 _19266_/D sky130_fd_sc_hd__o21a_1
XFILLER_235_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13953_ _13945_/B2 _13942_/X _13944_/Y _13952_/Y vssd1 vssd1 vccd1 vccd1 _14036_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_143_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19460_ _19526_/CLK _19460_/D vssd1 vssd1 vccd1 vccd1 _19460_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12904_ _09866_/Y _13292_/A2 _12903_/X _13256_/B1 _17922_/Q vssd1 vssd1 vccd1 vccd1
+ _12905_/B sky130_fd_sc_hd__a32o_1
X_16672_ _19245_/Q _16674_/C _16671_/Y vssd1 vssd1 vccd1 vccd1 _19245_/D sky130_fd_sc_hd__o21a_1
XFILLER_207_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13884_ _19389_/Q _13884_/A2 _13882_/X _13883_/X _13884_/C1 vssd1 vssd1 vccd1 vccd1
+ _13884_/X sky130_fd_sc_hd__o221a_4
XFILLER_185_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18411_ _19592_/CLK _18411_/D vssd1 vssd1 vccd1 vccd1 _18411_/Q sky130_fd_sc_hd__dfxtp_1
X_15623_ _15623_/A _15662_/C _15623_/C vssd1 vssd1 vccd1 vccd1 _15625_/B sky130_fd_sc_hd__or3_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ _19553_/CLK _19391_/D vssd1 vssd1 vccd1 vccd1 _19391_/Q sky130_fd_sc_hd__dfxtp_1
X_12835_ _12835_/A _12835_/B vssd1 vssd1 vccd1 vccd1 _12835_/Y sky130_fd_sc_hd__nor2_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _19620_/CLK _18342_/D vssd1 vssd1 vccd1 vccd1 _18342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15554_/A _15554_/B vssd1 vssd1 vccd1 vccd1 _15557_/C sky130_fd_sc_hd__or2_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12766_/A0 _09980_/Y _13446_/B vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _17707_/A0 _18355_/Q _14521_/S vssd1 vssd1 vccd1 vccd1 _18355_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11717_ _18531_/Q _18530_/Q vssd1 vssd1 vccd1 vccd1 _14417_/C sky130_fd_sc_hd__nand2b_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _19640_/CLK _18273_/D vssd1 vssd1 vccd1 vccd1 _18273_/Q sky130_fd_sc_hd__dfxtp_4
X_12697_ _12614_/B _12648_/B _12729_/B vssd1 vssd1 vccd1 vccd1 _12697_/X sky130_fd_sc_hd__mux2_1
X_15485_ _15508_/B vssd1 vssd1 vccd1 vccd1 _15485_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17224_ _18102_/Q _17382_/A _17123_/Y _17241_/B vssd1 vssd1 vccd1 vccd1 _17224_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14436_ _18575_/Q _14450_/B vssd1 vssd1 vccd1 vccd1 _18288_/D sky130_fd_sc_hd__and2_1
X_11648_ _12603_/B _12796_/S vssd1 vssd1 vccd1 vccd1 _11650_/B sky130_fd_sc_hd__and2b_1
XFILLER_122_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 core_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_2
Xinput23 core_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput34 core_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17155_ _19403_/Q _17124_/B _17448_/A _17212_/B2 vssd1 vssd1 vccd1 vccd1 _17156_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xinput45 dout0[11] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11579_ _11579_/A _11579_/B vssd1 vssd1 vccd1 vccd1 _11579_/Y sky130_fd_sc_hd__nor2_1
X_14367_ _18219_/Q _17674_/A0 _14377_/S vssd1 vssd1 vccd1 vccd1 _18219_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput56 dout0[21] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput67 dout0[31] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_2
X_16106_ _16140_/A1 _16105_/Y _16149_/A vssd1 vssd1 vccd1 vccd1 _18755_/D sky130_fd_sc_hd__a21oi_1
Xinput78 dout0[41] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput89 dout0[51] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_2
X_13318_ _14154_/B1 _13313_/X _13317_/X _11523_/B _12442_/C vssd1 vssd1 vccd1 vccd1
+ _13318_/X sky130_fd_sc_hd__o221a_1
XFILLER_182_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14298_ _17716_/A0 _18157_/Q _14305_/S vssd1 vssd1 vccd1 vccd1 _18157_/D sky130_fd_sc_hd__mux2_1
X_17086_ _17169_/B _17108_/A2 _17085_/X _17360_/A vssd1 vssd1 vccd1 vccd1 _19376_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16037_ _16038_/A _18732_/Q _16046_/A _16036_/Y vssd1 vssd1 vccd1 vccd1 _18731_/D
+ sky130_fd_sc_hd__o211a_1
X_13249_ _17865_/Q _13945_/A2 _13241_/X _13945_/B2 _13952_/B1 vssd1 vssd1 vccd1 vccd1
+ _13249_/X sky130_fd_sc_hd__a221o_1
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17988_ _19622_/CLK _17988_/D vssd1 vssd1 vccd1 vccd1 _17988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16939_ _19319_/Q _17190_/B _16947_/S vssd1 vssd1 vccd1 vccd1 _16940_/B sky130_fd_sc_hd__mux2_1
Xfanout1880 _17330_/A vssd1 vssd1 vccd1 vccd1 _17159_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_266_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1891 _16110_/B1 vssd1 vssd1 vccd1 vccd1 _16128_/B1 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_146_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19507_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09411_ _09718_/S _09406_/X _09410_/X vssd1 vssd1 vccd1 vccd1 _09411_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_252_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18609_ _19589_/CLK _18609_/D vssd1 vssd1 vccd1 vccd1 _18609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19589_ _19589_/CLK _19589_/D vssd1 vssd1 vccd1 vccd1 _19589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09342_ _19043_/Q _19011_/Q _10099_/S vssd1 vssd1 vccd1 vccd1 _09342_/X sky130_fd_sc_hd__mux2_1
XFILLER_279_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09273_ _10409_/A _09271_/X _09272_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09274_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_221_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08988_ input126/X input161/X _09657_/S vssd1 vssd1 vccd1 vccd1 _08988_/X sky130_fd_sc_hd__mux2_8
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10950_ _12320_/B _11135_/S _11181_/B1 _10949_/Y vssd1 vssd1 vccd1 vccd1 _10985_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09609_ _11210_/A1 _09611_/B _09608_/Y _11055_/B2 vssd1 vssd1 vccd1 vccd1 _15194_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_244_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10881_ _18646_/Q _18068_/Q _19087_/Q _18991_/Q _10500_/S _10881_/S1 vssd1 vssd1
+ vccd1 vccd1 _10882_/B sky130_fd_sc_hd__mux4_1
XFILLER_244_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12620_ _13188_/B _13188_/C _13188_/A vssd1 vssd1 vccd1 vccd1 _13225_/C sky130_fd_sc_hd__o21a_1
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12551_ _12552_/A _12552_/B vssd1 vssd1 vccd1 vccd1 _12551_/Y sky130_fd_sc_hd__nor2_2
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11502_ _09374_/S _11499_/X _11501_/X vssd1 vssd1 vccd1 vccd1 _11502_/Y sky130_fd_sc_hd__a21oi_4
XPHY_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12482_ _17919_/Q _12285_/A _12482_/S vssd1 vssd1 vccd1 vccd1 _12553_/A sky130_fd_sc_hd__mux2_2
X_15270_ _18570_/Q _18569_/Q _15270_/C vssd1 vssd1 vccd1 vccd1 _15314_/C sky130_fd_sc_hd__and3_2
XFILLER_184_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11433_ _11511_/A _11433_/B vssd1 vssd1 vccd1 vccd1 _11433_/Y sky130_fd_sc_hd__nand2_1
XFILLER_200_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14221_ _18282_/Q _14224_/B _14220_/Y _14430_/B vssd1 vssd1 vccd1 vccd1 _18108_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14152_ _14152_/A _14152_/B _14152_/C vssd1 vssd1 vccd1 vccd1 _14153_/D sky130_fd_sc_hd__nor3_4
XFILLER_165_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11364_ _11131_/A _11343_/Y _11349_/Y _11356_/Y _11363_/X vssd1 vssd1 vccd1 vccd1
+ _11364_/X sky130_fd_sc_hd__o32a_4
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13103_ _15911_/A _12536_/Y _12505_/Y vssd1 vssd1 vccd1 vccd1 _13103_/X sky130_fd_sc_hd__a21o_1
XFILLER_217_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10315_ _10313_/X _10314_/X _10315_/S vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14083_ _16500_/A0 _18023_/Q _14104_/S vssd1 vssd1 vccd1 vccd1 _18023_/D sky130_fd_sc_hd__mux2_1
X_18960_ _19226_/CLK _18960_/D vssd1 vssd1 vccd1 vccd1 _18960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11295_ _17966_/Q _11295_/A2 _11371_/B1 vssd1 vssd1 vccd1 vccd1 _11295_/X sky130_fd_sc_hd__a21o_1
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17911_ _18817_/CLK _17911_/D vssd1 vssd1 vccd1 vccd1 _17911_/Q sky130_fd_sc_hd__dfxtp_1
X_13034_ _13032_/Y _13083_/C vssd1 vssd1 vccd1 vccd1 _14142_/B sky130_fd_sc_hd__and2b_1
XFILLER_279_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10246_ _10253_/A _10245_/X _10244_/X vssd1 vssd1 vccd1 vccd1 _10246_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18891_ _19622_/CLK _18891_/D vssd1 vssd1 vccd1 vccd1 _18891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1110 _12586_/X vssd1 vssd1 vccd1 vccd1 _13758_/A sky130_fd_sc_hd__buf_6
XFILLER_105_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1121 _12437_/Y vssd1 vssd1 vccd1 vccd1 _13289_/A sky130_fd_sc_hd__buf_4
X_17842_ _19363_/CLK _17842_/D vssd1 vssd1 vccd1 vccd1 _17842_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1132 _13970_/B2 vssd1 vssd1 vccd1 vccd1 _13869_/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_239_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10177_ _11017_/A1 _18162_/Q _18808_/Q _10176_/S vssd1 vssd1 vccd1 vccd1 _10177_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_267_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1143 _10194_/C1 vssd1 vssd1 vccd1 vccd1 _09859_/A sky130_fd_sc_hd__buf_8
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1154 _09083_/A vssd1 vssd1 vccd1 vccd1 _15120_/A sky130_fd_sc_hd__buf_6
Xfanout1165 _15948_/B1 vssd1 vssd1 vccd1 vccd1 _15923_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1176 _14204_/S vssd1 vssd1 vccd1 vccd1 _14200_/S sky130_fd_sc_hd__buf_6
XFILLER_248_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17773_ _19601_/CLK _17773_/D vssd1 vssd1 vccd1 vccd1 _17773_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1187 _10083_/X vssd1 vssd1 vccd1 vccd1 _11064_/B1 sky130_fd_sc_hd__clkbuf_2
X_14985_ _18130_/Q _14671_/X _14934_/X _14984_/X vssd1 vssd1 vccd1 vccd1 _14985_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1198 _13797_/A0 vssd1 vssd1 vccd1 vccd1 _14155_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_281_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19512_ _19546_/CLK _19512_/D vssd1 vssd1 vccd1 vccd1 _19512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16724_ _16795_/A _16724_/B _16729_/C vssd1 vssd1 vccd1 vccd1 _19260_/D sky130_fd_sc_hd__nor3_1
XFILLER_263_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13936_ _15382_/B2 _13932_/X _13935_/Y _13936_/B2 vssd1 vssd1 vccd1 vccd1 _13937_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_240_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19443_ _19444_/CLK _19443_/D vssd1 vssd1 vccd1 vccd1 _19443_/Q sky130_fd_sc_hd__dfxtp_1
X_16655_ _16768_/A _16661_/C vssd1 vssd1 vccd1 vccd1 _16655_/Y sky130_fd_sc_hd__nor2_1
XFILLER_263_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13867_ _13323_/B _13865_/X _13866_/X _13968_/A1 vssd1 vssd1 vccd1 vccd1 _13867_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_234_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15606_ _15623_/A _15602_/Y _15605_/X vssd1 vssd1 vccd1 vccd1 _15606_/X sky130_fd_sc_hd__a21o_1
X_19374_ _19458_/CLK _19374_/D vssd1 vssd1 vccd1 vccd1 _19374_/Q sky130_fd_sc_hd__dfxtp_1
X_12818_ _12714_/X _12730_/Y _12818_/S vssd1 vssd1 vccd1 vccd1 _12818_/X sky130_fd_sc_hd__mux2_1
X_16586_ _16619_/A0 _19190_/Q _16586_/S vssd1 vssd1 vccd1 vccd1 _19190_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13798_ _13962_/B _13797_/X _10454_/B vssd1 vssd1 vccd1 vccd1 _13798_/X sky130_fd_sc_hd__a21o_1
X_18325_ _19604_/CLK _18325_/D vssd1 vssd1 vccd1 vccd1 _18325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ _15789_/A1 _15536_/Y _15537_/B1 vssd1 vssd1 vccd1 vccd1 _15538_/C sky130_fd_sc_hd__a21oi_1
XFILLER_176_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12749_ _12746_/B _12748_/Y _12935_/S vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18256_ _19638_/CLK _18256_/D vssd1 vssd1 vccd1 vccd1 _18256_/Q sky130_fd_sc_hd__dfxtp_1
X_15468_ _19440_/Q _15124_/B _15731_/B1 _15467_/X vssd1 vssd1 vccd1 vccd1 _15468_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17207_ _17210_/A _17207_/B vssd1 vssd1 vccd1 vccd1 _19420_/D sky130_fd_sc_hd__nor2_1
X_14419_ _19228_/Q _15014_/B _18274_/D vssd1 vssd1 vccd1 vccd1 _18270_/D sky130_fd_sc_hd__and3_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18187_ _19146_/CLK _18187_/D vssd1 vssd1 vccd1 vccd1 _18187_/Q sky130_fd_sc_hd__dfxtp_1
X_15399_ _15399_/A _15399_/B vssd1 vssd1 vccd1 vccd1 _15399_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_265_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17138_ _17141_/A _17138_/B vssd1 vssd1 vccd1 vccd1 _19397_/D sky130_fd_sc_hd__nor2_1
XFILLER_171_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09960_ _18440_/Q _18341_/Q _10281_/S vssd1 vssd1 vccd1 vccd1 _09960_/X sky130_fd_sc_hd__mux2_1
X_17069_ _19368_/Q _17077_/B vssd1 vssd1 vccd1 vccd1 _17069_/X sky130_fd_sc_hd__or2_1
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08911_ _08932_/A _17795_/Q vssd1 vssd1 vccd1 vccd1 _08942_/B sky130_fd_sc_hd__nand2b_2
XFILLER_131_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _11274_/S1 _09880_/X _09890_/X _08950_/A vssd1 vssd1 vccd1 vccd1 _09891_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08842_ _09690_/A vssd1 vssd1 vccd1 vccd1 _08842_/Y sky130_fd_sc_hd__clkinv_2
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09325_ _11217_/A _09902_/B _09325_/C _09325_/D vssd1 vssd1 vccd1 vccd1 _09326_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_159_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ _19044_/Q _19012_/Q _11481_/C vssd1 vssd1 vccd1 vccd1 _09256_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19645_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09187_ _11484_/B1 _09178_/X _11466_/B1 vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__a21o_1
XFILLER_181_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10100_ _10098_/X _10099_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _10100_/X sky130_fd_sc_hd__mux2_2
XFILLER_255_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11080_ _11305_/A1 _17775_/Q _11309_/S _18324_/Q _10784_/S vssd1 vssd1 vccd1 vccd1
+ _11080_/X sky130_fd_sc_hd__o221a_1
XFILLER_122_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput202 localMemory_wb_adr_i[20] vssd1 vssd1 vccd1 vccd1 _12269_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10031_ _18236_/Q _18811_/Q _10500_/S vssd1 vssd1 vccd1 vccd1 _10031_/X sky130_fd_sc_hd__mux2_1
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput213 localMemory_wb_adr_i[9] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__clkbuf_2
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput224 localMemory_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input224/X sky130_fd_sc_hd__buf_8
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput235 localMemory_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 input235/X sky130_fd_sc_hd__buf_12
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput246 localMemory_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input246/X sky130_fd_sc_hd__buf_8
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput257 manufacturerID[3] vssd1 vssd1 vccd1 vccd1 _15866_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput268 partID[13] vssd1 vssd1 vccd1 vccd1 input268/X sky130_fd_sc_hd__clkbuf_2
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput279 partID[9] vssd1 vssd1 vccd1 vccd1 _15917_/A sky130_fd_sc_hd__buf_2
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14770_ _14768_/X _14769_/X _14913_/B1 vssd1 vssd1 vccd1 vccd1 _14770_/X sky130_fd_sc_hd__a21o_1
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _16054_/A _16034_/S _16069_/B vssd1 vssd1 vccd1 vccd1 _15849_/A sky130_fd_sc_hd__nor3_4
XFILLER_216_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13721_ _19384_/Q _13884_/A2 _13719_/X _13720_/X _13884_/C1 vssd1 vssd1 vccd1 vccd1
+ _13721_/X sky130_fd_sc_hd__o221a_4
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10933_ _11327_/S _11572_/A1 _19214_/Q _11578_/S vssd1 vssd1 vccd1 vccd1 _10933_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_244_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16440_ _19048_/Q _11376_/B _16454_/S vssd1 vssd1 vccd1 vccd1 _19048_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10864_ _18863_/Q _18895_/Q _10864_/S vssd1 vssd1 vccd1 vccd1 _10864_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13652_ _19544_/Q _13921_/S vssd1 vssd1 vccd1 vccd1 _13652_/X sky130_fd_sc_hd__or2_1
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ _12796_/S _12603_/B vssd1 vssd1 vccd1 vccd1 _12842_/B sky130_fd_sc_hd__or2_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _16471_/A0 _18982_/Q _16390_/S vssd1 vssd1 vccd1 vccd1 _18982_/D sky130_fd_sc_hd__mux2_1
XFILLER_223_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _17843_/Q _13846_/B _12548_/X vssd1 vssd1 vccd1 vccd1 _13583_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_169_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10795_ _18328_/Q _17779_/Q _11604_/S vssd1 vssd1 vccd1 vccd1 _10795_/X sky130_fd_sc_hd__mux2_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18110_ _18778_/CLK _18110_/D vssd1 vssd1 vccd1 vccd1 _18110_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_158_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _19465_/Q _19399_/Q _15299_/B vssd1 vssd1 vccd1 vccd1 _15322_/X sky130_fd_sc_hd__a21o_1
X_12534_ _19296_/Q _13174_/A _12533_/Y input1/X _12531_/X vssd1 vssd1 vccd1 vccd1
+ _12534_/X sky130_fd_sc_hd__a221o_4
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _19154_/CLK _19090_/D vssd1 vssd1 vccd1 vccd1 _19090_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18041_ _19611_/CLK _18041_/D vssd1 vssd1 vccd1 vccd1 _18041_/Q sky130_fd_sc_hd__dfxtp_1
X_15253_ _15228_/Y _15233_/B _15230_/B vssd1 vssd1 vccd1 vccd1 _15254_/B sky130_fd_sc_hd__o21ai_4
X_12465_ _16852_/A _09777_/A _16839_/A vssd1 vssd1 vccd1 vccd1 _12499_/A sky130_fd_sc_hd__a21bo_2
X_14204_ _18713_/Q _18100_/Q _14204_/S vssd1 vssd1 vccd1 vccd1 _14205_/B sky130_fd_sc_hd__mux2_1
X_11416_ _11414_/X _11415_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _11416_/X sky130_fd_sc_hd__mux2_1
X_12396_ _12429_/A1 _12409_/A2 _09035_/X _12417_/B1 _18392_/Q vssd1 vssd1 vccd1 vccd1
+ _12397_/B sky130_fd_sc_hd__o32ai_2
X_15184_ _19428_/Q _15140_/B _15731_/B1 _15183_/X vssd1 vssd1 vccd1 vccd1 _15192_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_153_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14135_ _16486_/A0 _18074_/Q _14137_/S vssd1 vssd1 vccd1 vccd1 _18074_/D sky130_fd_sc_hd__mux2_1
X_11347_ _18857_/Q _18889_/Q _19049_/Q _19017_/Q _11360_/B2 _11357_/S1 vssd1 vssd1
+ vccd1 vccd1 _11347_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18943_ _19592_/CLK _18943_/D vssd1 vssd1 vccd1 vccd1 _18943_/Q sky130_fd_sc_hd__dfxtp_1
X_14066_ _17683_/A0 _18008_/Q _14073_/S vssd1 vssd1 vccd1 vccd1 _18008_/D sky130_fd_sc_hd__mux2_1
X_11278_ _11276_/X _11277_/X _11285_/S vssd1 vssd1 vccd1 vccd1 _11278_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10229_ _11210_/A1 _10166_/X _10228_/X _09523_/A vssd1 vssd1 vccd1 vccd1 _13874_/A
+ sky130_fd_sc_hd__a22o_4
X_13017_ _19429_/Q _12560_/B _13015_/X _13016_/X _12560_/A vssd1 vssd1 vccd1 vccd1
+ _13017_/X sky130_fd_sc_hd__o221a_1
X_18874_ _19055_/CLK _18874_/D vssd1 vssd1 vccd1 vccd1 _18874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17825_ _18713_/CLK _17825_/D vssd1 vssd1 vccd1 vccd1 _17825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17756_ _18656_/Q vssd1 vssd1 vccd1 vccd1 _18656_/D sky130_fd_sc_hd__clkbuf_2
X_14968_ _14968_/A vssd1 vssd1 vccd1 vccd1 _14968_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_94_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16707_ _16795_/A _16713_/C vssd1 vssd1 vccd1 vccd1 _16707_/Y sky130_fd_sc_hd__nor2_1
XFILLER_223_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13919_ _19262_/Q _13943_/A2 _13943_/B1 _19294_/Q vssd1 vssd1 vccd1 vccd1 _13919_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17687_ _17720_/A0 _19614_/Q _17687_/S vssd1 vssd1 vccd1 vccd1 _19614_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14899_ _14895_/X _14898_/X _15010_/B1 vssd1 vssd1 vccd1 vccd1 _14899_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19426_ _19492_/CLK _19426_/D vssd1 vssd1 vccd1 vccd1 _19426_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16638_ _19235_/Q _19234_/Q _16677_/A vssd1 vssd1 vccd1 vccd1 _16643_/C sky130_fd_sc_hd__and3_1
XFILLER_222_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19357_ _19485_/CLK _19357_/D vssd1 vssd1 vccd1 vccd1 _19357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16569_ _16602_/A0 _19173_/Q _16589_/S vssd1 vssd1 vccd1 vccd1 _19173_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09110_ _09457_/B _18886_/Q _09285_/C vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__and3_1
X_18308_ _19047_/CLK _18308_/D vssd1 vssd1 vccd1 vccd1 _18308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19288_ _19291_/CLK _19288_/D vssd1 vssd1 vccd1 vccd1 _19288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ _09042_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _11687_/A sky130_fd_sc_hd__and2_4
XFILLER_198_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18239_ _19621_/CLK _18239_/D vssd1 vssd1 vccd1 vccd1 _18239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09943_ _17896_/Q _15120_/A vssd1 vssd1 vccd1 vccd1 _09943_/Y sky130_fd_sc_hd__nor2_1
Xfanout903 _09248_/X vssd1 vssd1 vccd1 vccd1 _16204_/A0 sky130_fd_sc_hd__buf_6
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout914 _16388_/S vssd1 vssd1 vccd1 vccd1 _16390_/S sky130_fd_sc_hd__buf_12
XFILLER_225_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout925 _16222_/S vssd1 vssd1 vccd1 vccd1 _16225_/S sky130_fd_sc_hd__clkbuf_16
Xfanout936 _14982_/B vssd1 vssd1 vccd1 vccd1 _15002_/B sky130_fd_sc_hd__clkbuf_4
Xfanout947 _14670_/Y vssd1 vssd1 vccd1 vccd1 _14964_/B1 sky130_fd_sc_hd__buf_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_161_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19506_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09874_ _08901_/A _18596_/Q _18167_/Q _10054_/S _08874_/D vssd1 vssd1 vccd1 vccd1
+ _09874_/X sky130_fd_sc_hd__a221o_1
Xfanout958 _14517_/S vssd1 vssd1 vccd1 vccd1 _14520_/S sky130_fd_sc_hd__buf_12
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout969 _14041_/Y vssd1 vssd1 vccd1 vccd1 _14073_/S sky130_fd_sc_hd__buf_12
XFILLER_285_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08825_ _08825_/A vssd1 vssd1 vccd1 vccd1 _15845_/A sky130_fd_sc_hd__inv_4
XFILLER_246_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_307 _18113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_318 _18104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_329 _11899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09308_ _09967_/S _09306_/X _09307_/X _11507_/S vssd1 vssd1 vccd1 vccd1 _09308_/X
+ sky130_fd_sc_hd__a211o_1
X_10580_ _11131_/A _10574_/X _10577_/X _10579_/X vssd1 vssd1 vccd1 vccd1 _10580_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09239_ _09033_/X _09238_/Y _09326_/A vssd1 vssd1 vccd1 vccd1 _09239_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _17883_/Q _12253_/C vssd1 vssd1 vccd1 vccd1 _12251_/B sky130_fd_sc_hd__and2_1
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11201_ _10371_/S _11198_/X _11200_/X vssd1 vssd1 vccd1 vccd1 _11201_/X sky130_fd_sc_hd__a21o_1
X_12181_ _17857_/Q _12184_/C _12187_/A vssd1 vssd1 vccd1 vccd1 _12181_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_269_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11132_ _11117_/Y _11130_/X _11131_/X vssd1 vssd1 vccd1 vccd1 _11132_/X sky130_fd_sc_hd__o21a_2
XFILLER_134_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15940_ _18689_/Q _15946_/A2 _15939_/X _15946_/C1 vssd1 vssd1 vccd1 vccd1 _18689_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ _12593_/A vssd1 vssd1 vccd1 vccd1 _13533_/A sky130_fd_sc_hd__inv_2
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ _18439_/Q _18340_/Q _11070_/S vssd1 vssd1 vccd1 vccd1 _10014_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_264_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15871_ _18666_/Q _15949_/A2 _15869_/X _15870_/X _15910_/C1 vssd1 vssd1 vccd1 vccd1
+ _18666_/D sky130_fd_sc_hd__o221a_1
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _19546_/Q _17622_/A2 _17591_/X _17193_/B _17609_/X vssd1 vssd1 vccd1 vccd1
+ _19546_/D sky130_fd_sc_hd__o221a_1
XFILLER_64_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ _14995_/A1 _14820_/X _14821_/X _14771_/X vssd1 vssd1 vccd1 vccd1 _14822_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _19453_/CLK _18590_/D vssd1 vssd1 vccd1 vccd1 _18590_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17541_ _17208_/Y _17493_/B _17540_/Y _16048_/A vssd1 vssd1 vccd1 vccd1 _17541_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_233_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _18107_/Q _14801_/B _14690_/Y _14752_/X vssd1 vssd1 vccd1 vccd1 _14753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _18511_/Q _11720_/X _11915_/X _11968_/B2 vssd1 vssd1 vccd1 vccd1 _11965_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _18124_/Q _18123_/Q _13704_/C vssd1 vssd1 vccd1 vccd1 _13736_/B sky130_fd_sc_hd__and3_1
XFILLER_233_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17472_ _18117_/Q _17539_/C1 _17470_/X _17471_/X vssd1 vssd1 vccd1 vccd1 _17472_/X
+ sky130_fd_sc_hd__a22o_1
X_10916_ _18645_/Q _18067_/Q _11581_/S vssd1 vssd1 vccd1 vccd1 _10916_/X sky130_fd_sc_hd__mux2_1
X_14684_ _14674_/X _14678_/X _14714_/B vssd1 vssd1 vccd1 vccd1 _14684_/X sky130_fd_sc_hd__a21o_1
XFILLER_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11896_ _11896_/A _11901_/B vssd1 vssd1 vccd1 vccd1 _11896_/X sky130_fd_sc_hd__or2_1
X_19211_ _19211_/CLK _19211_/D vssd1 vssd1 vccd1 vccd1 _19211_/Q sky130_fd_sc_hd__dfxtp_1
X_16423_ _16621_/A0 _19032_/Q _16424_/S vssd1 vssd1 vccd1 vccd1 _19032_/D sky130_fd_sc_hd__mux2_1
XFILLER_260_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13635_ _13682_/B2 _13624_/X _13626_/Y _13634_/Y vssd1 vssd1 vccd1 vccd1 _14016_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10847_ _18036_/Q _18004_/Q _10853_/S vssd1 vssd1 vccd1 vccd1 _10847_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19142_ _19142_/CLK _19142_/D vssd1 vssd1 vccd1 vccd1 _19142_/Q sky130_fd_sc_hd__dfxtp_1
X_16354_ _18966_/Q _16553_/A0 _16357_/S vssd1 vssd1 vccd1 vccd1 _18966_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13566_ _13566_/A _13961_/A vssd1 vssd1 vccd1 vccd1 _13566_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ _11572_/A1 _17779_/Q _10853_/S _18328_/Q vssd1 vssd1 vccd1 vccd1 _10778_/X
+ sky130_fd_sc_hd__o22a_1
X_15305_ _18111_/Q _15133_/Y _15304_/X _15382_/B2 vssd1 vssd1 vccd1 vccd1 _15305_/X
+ sky130_fd_sc_hd__a22o_1
X_12517_ _12768_/A _12584_/A vssd1 vssd1 vccd1 vccd1 _13925_/S sky130_fd_sc_hd__or2_4
X_19073_ _19147_/CLK _19073_/D vssd1 vssd1 vccd1 vccd1 _19073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16285_ _16418_/A0 _18899_/Q _16292_/S vssd1 vssd1 vccd1 vccd1 _18899_/D sky130_fd_sc_hd__mux2_1
XFILLER_200_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13497_ _19539_/Q _13921_/S vssd1 vssd1 vccd1 vccd1 _13497_/X sky130_fd_sc_hd__or2_1
XFILLER_172_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18024_ _19213_/CLK _18024_/D vssd1 vssd1 vccd1 vccd1 _18024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15236_ _17382_/A _15236_/B _15236_/C vssd1 vssd1 vccd1 vccd1 _15236_/Y sky130_fd_sc_hd__nor3_1
XFILLER_161_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ _13185_/A _12761_/B _12448_/C _12448_/D vssd1 vssd1 vccd1 vccd1 _15083_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_172_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ _15167_/A _15167_/B vssd1 vssd1 vccd1 vccd1 _15167_/Y sky130_fd_sc_hd__xnor2_1
X_12379_ _12379_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14118_ _16535_/A0 _18057_/Q _14139_/S vssd1 vssd1 vccd1 vccd1 _18057_/D sky130_fd_sc_hd__mux2_1
XFILLER_153_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098_ _19377_/Q _15086_/B input178/X _15097_/X vssd1 vssd1 vccd1 vccd1 _15101_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14049_ _17666_/A0 _17991_/Q _14070_/S vssd1 vssd1 vccd1 vccd1 _17991_/D sky130_fd_sc_hd__mux2_1
X_18926_ _19637_/CLK _18926_/D vssd1 vssd1 vccd1 vccd1 _18926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18857_ _19216_/CLK _18857_/D vssd1 vssd1 vccd1 vccd1 _18857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09590_ _09588_/X _09589_/X _10371_/S vssd1 vssd1 vccd1 vccd1 _09590_/X sky130_fd_sc_hd__mux2_1
X_17808_ _17814_/CLK _17808_/D vssd1 vssd1 vccd1 vccd1 _17808_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_269_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18788_ _19627_/CLK _18788_/D vssd1 vssd1 vccd1 vccd1 _18788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17739_ _18639_/Q vssd1 vssd1 vccd1 vccd1 _18639_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_270_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19409_ _19507_/CLK _19409_/D vssd1 vssd1 vccd1 vccd1 _19409_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09024_ _09021_/X _09022_/X _09023_/X _08927_/Y vssd1 vssd1 vccd1 vccd1 _09025_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_148_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout700 _12545_/Y vssd1 vssd1 vccd1 vccd1 _13425_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout711 _13115_/C1 vssd1 vssd1 vccd1 vccd1 _13952_/B1 sky130_fd_sc_hd__buf_6
Xfanout1709 _12488_/B vssd1 vssd1 vccd1 vccd1 _09750_/S sky130_fd_sc_hd__buf_8
XFILLER_132_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout722 _12497_/Y vssd1 vssd1 vccd1 vccd1 _13942_/B1 sky130_fd_sc_hd__buf_6
X_09926_ _10262_/A1 _18595_/Q _18166_/Q _09671_/S _10315_/S vssd1 vssd1 vccd1 vccd1
+ _09926_/X sky130_fd_sc_hd__a221o_1
Xfanout733 _16539_/A0 vssd1 vssd1 vccd1 vccd1 _17672_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_131_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout744 _12878_/S vssd1 vssd1 vccd1 vccd1 _12942_/S sky130_fd_sc_hd__buf_4
XFILLER_86_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout755 _12739_/S vssd1 vssd1 vccd1 vccd1 _13136_/S sky130_fd_sc_hd__buf_6
XFILLER_274_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout766 _17723_/S vssd1 vssd1 vccd1 vccd1 _17719_/S sky130_fd_sc_hd__buf_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09857_ _09857_/A1 _09853_/X _09856_/X _11237_/B1 vssd1 vssd1 vccd1 vccd1 _09857_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout777 _16623_/S vssd1 vssd1 vccd1 vccd1 _16618_/S sky130_fd_sc_hd__buf_12
Xfanout788 _16525_/Y vssd1 vssd1 vccd1 vccd1 _16554_/S sky130_fd_sc_hd__clkbuf_16
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout799 _16325_/S vssd1 vssd1 vccd1 vccd1 _16324_/S sky130_fd_sc_hd__clkbuf_16
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09788_ _09784_/X _09785_/X _10040_/S vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__mux2_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_104 _13941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_115 _11846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_137 _11836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _11868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11750_/A _11750_/B vssd1 vssd1 vccd1 vccd1 _11751_/A sky130_fd_sc_hd__xnor2_4
XFILLER_242_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_159 _11972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10701_ _10699_/X _10700_/X _10706_/S vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__mux2_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11681_ _11681_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _13330_/B sky130_fd_sc_hd__xnor2_4
XFILLER_186_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13420_ _13409_/Y _13412_/Y _13419_/X _13966_/C1 vssd1 vssd1 vccd1 vccd1 _13420_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10632_ _10630_/X _10631_/X _10632_/S vssd1 vssd1 vccd1 vccd1 _10633_/B sky130_fd_sc_hd__mux2_1
XFILLER_197_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10563_ _10532_/A _10562_/X _10532_/Y _11790_/B vssd1 vssd1 vccd1 vccd1 _10564_/B
+ sky130_fd_sc_hd__a211o_1
X_13351_ _13351_/A _13351_/B vssd1 vssd1 vccd1 vccd1 _14145_/A sky130_fd_sc_hd__xor2_1
XFILLER_210_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _14417_/C _12271_/B _12276_/B _15835_/C vssd1 vssd1 vccd1 vccd1 _16819_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_10_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16070_ _16054_/A _16063_/B _08825_/A vssd1 vssd1 vccd1 vccd1 _16070_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13282_ _15923_/A _12575_/Y _13276_/X _13427_/A1 vssd1 vssd1 vccd1 vccd1 _13282_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _10817_/A1 _19579_/Q _10500_/S _19611_/Q _10033_/S vssd1 vssd1 vccd1 vccd1
+ _10494_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15021_ _18510_/Q input210/X _15024_/S vssd1 vssd1 vccd1 vccd1 _18510_/D sky130_fd_sc_hd__mux2_1
X_12233_ _12241_/A _12233_/B _12234_/B vssd1 vssd1 vccd1 vccd1 _17876_/D sky130_fd_sc_hd__nor3_1
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ _17850_/Q _12162_/B _12163_/Y vssd1 vssd1 vccd1 vccd1 _17850_/D sky130_fd_sc_hd__o21a_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _11113_/X _11114_/X _11127_/S vssd1 vssd1 vccd1 vccd1 _11115_/X sky130_fd_sc_hd__mux2_1
X_12095_ _17823_/Q _17824_/Q _17825_/Q vssd1 vssd1 vccd1 vccd1 _12100_/C sky130_fd_sc_hd__and3_2
X_16972_ _16972_/A _16972_/B vssd1 vssd1 vccd1 vccd1 _19327_/D sky130_fd_sc_hd__and2_1
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15923_ _15923_/A _15941_/S _15923_/C vssd1 vssd1 vccd1 vccd1 _15923_/X sky130_fd_sc_hd__and3_1
X_11046_ _18550_/Q _18425_/Q _18034_/Q _18002_/Q _11426_/B2 _11046_/S1 vssd1 vssd1
+ vccd1 vccd1 _11046_/X sky130_fd_sc_hd__mux4_1
X_18711_ _18713_/CLK _18711_/D vssd1 vssd1 vccd1 vccd1 _18711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18642_ _19133_/CLK _18642_/D vssd1 vssd1 vccd1 vccd1 _18642_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _15854_/A _15854_/B vssd1 vssd1 vccd1 vccd1 _15854_/Y sky130_fd_sc_hd__nand2_1
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _14805_/A vssd1 vssd1 vccd1 vccd1 _14805_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18573_ _19433_/CLK _18573_/D vssd1 vssd1 vccd1 vccd1 _18573_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_224_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _13941_/A _15502_/B _13969_/Y _15112_/B vssd1 vssd1 vccd1 vccd1 _15785_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12997_ _12997_/A vssd1 vssd1 vccd1 vccd1 _12997_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _17390_/Y _17521_/X _17522_/X _17523_/X _17380_/A vssd1 vssd1 vccd1 vccd1
+ _19516_/D sky130_fd_sc_hd__o311a_1
XFILLER_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _14865_/A1 _14735_/X _14865_/B1 vssd1 vssd1 vccd1 vccd1 _14736_/Y sky130_fd_sc_hd__o21ai_2
X_11948_ _11953_/B2 _11894_/B _11894_/C _11953_/A2 input235/X vssd1 vssd1 vccd1 vccd1
+ _11948_/X sky130_fd_sc_hd__a32o_4
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17455_ _13366_/B _15118_/A _15117_/A _17803_/Q _15116_/B vssd1 vssd1 vccd1 vccd1
+ _17455_/X sky130_fd_sc_hd__a221o_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14667_ _14667_/A1 _14417_/B _15835_/A _14665_/X vssd1 vssd1 vccd1 vccd1 _14667_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_60_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11879_ _10489_/B _11864_/B _11926_/A1 vssd1 vssd1 vccd1 vccd1 _11882_/B sky130_fd_sc_hd__o21ai_2
X_16406_ _11452_/B _19015_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _19015_/D sky130_fd_sc_hd__mux2_1
X_13618_ _10831_/A _13912_/B1 _13912_/A2 _11537_/B _14153_/A vssd1 vssd1 vccd1 vccd1
+ _13618_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17386_ _19489_/Q _17386_/B vssd1 vssd1 vccd1 vccd1 _17386_/X sky130_fd_sc_hd__and2_1
X_14598_ _14527_/B _14597_/X _14596_/A vssd1 vssd1 vccd1 vccd1 _18406_/D sky130_fd_sc_hd__o21ba_1
XFILLER_119_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19125_ _19157_/CLK _19125_/D vssd1 vssd1 vccd1 vccd1 _19125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16337_ _18949_/Q _17669_/A0 _16357_/S vssd1 vssd1 vccd1 vccd1 _18949_/D sky130_fd_sc_hd__mux2_1
X_13549_ _17842_/Q _13744_/A2 _13744_/B1 _17874_/Q vssd1 vssd1 vccd1 vccd1 _13549_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19056_ _19607_/CLK _19056_/D vssd1 vssd1 vccd1 vccd1 _19056_/Q sky130_fd_sc_hd__dfxtp_1
X_16268_ _17666_/A0 _18882_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _18882_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18007_ _19638_/CLK _18007_/D vssd1 vssd1 vccd1 vccd1 _18007_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput303 _19652_/X vssd1 vssd1 vccd1 vccd1 clk0 sky130_fd_sc_hd__clkbuf_2
X_15219_ _15219_/A _15219_/B vssd1 vssd1 vccd1 vccd1 _15263_/C sky130_fd_sc_hd__xnor2_4
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput314 _11762_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[18] sky130_fd_sc_hd__buf_4
X_16199_ _16431_/A1 _18815_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _18815_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput325 _11733_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[2] sky130_fd_sc_hd__buf_4
Xoutput336 _11818_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[11] sky130_fd_sc_hd__buf_4
XFILLER_114_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput347 _11863_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[21] sky130_fd_sc_hd__buf_4
Xoutput358 _11909_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[31] sky130_fd_sc_hd__buf_4
Xoutput369 _11781_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[3] sky130_fd_sc_hd__buf_4
XFILLER_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09711_ _18443_/Q _18344_/Q _09720_/S vssd1 vssd1 vccd1 vccd1 _09711_/X sky130_fd_sc_hd__mux2_1
XFILLER_256_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18909_ _19620_/CLK _18909_/D vssd1 vssd1 vccd1 vccd1 _18909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09642_ _09611_/A _09641_/X _09611_/Y _11790_/B vssd1 vssd1 vccd1 vccd1 _11796_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09573_ _09027_/A _09034_/B _09572_/X _10162_/B _09483_/Y vssd1 vssd1 vccd1 vccd1
+ _09574_/C sky130_fd_sc_hd__a32o_1
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09007_ _18268_/Q _18199_/Q vssd1 vssd1 vccd1 vccd1 _09007_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1506 fanout1514/X vssd1 vssd1 vccd1 vccd1 _10215_/S sky130_fd_sc_hd__buf_6
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1517 _09302_/S vssd1 vssd1 vccd1 vccd1 _09306_/S sky130_fd_sc_hd__buf_6
XFILLER_238_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout530 _11899_/A vssd1 vssd1 vccd1 vccd1 _11770_/B1 sky130_fd_sc_hd__buf_4
Xfanout1528 _10643_/S vssd1 vssd1 vccd1 vccd1 _11611_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_263_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1539 _09967_/S vssd1 vssd1 vccd1 vccd1 _10419_/S sky130_fd_sc_hd__buf_4
Xfanout541 _17540_/B1 vssd1 vssd1 vccd1 vccd1 _15782_/A1 sky130_fd_sc_hd__buf_4
X_09909_ _09028_/B _09908_/X _09042_/Y vssd1 vssd1 vccd1 vccd1 _09909_/Y sky130_fd_sc_hd__a21oi_1
Xfanout552 _15122_/Y vssd1 vssd1 vccd1 vccd1 _17202_/A sky130_fd_sc_hd__buf_8
Xfanout563 _15437_/B1 vssd1 vssd1 vccd1 vccd1 _15223_/A sky130_fd_sc_hd__buf_2
Xfanout574 _16096_/A1 vssd1 vssd1 vccd1 vccd1 _16142_/A1 sky130_fd_sc_hd__buf_4
XFILLER_219_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout585 _12024_/Y vssd1 vssd1 vccd1 vccd1 _12035_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12920_ _17826_/Q _12919_/X _13105_/B vssd1 vssd1 vccd1 vccd1 _12920_/X sky130_fd_sc_hd__mux2_2
Xfanout596 _14268_/B vssd1 vssd1 vccd1 vccd1 _14224_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_207_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _12851_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12851_/X sky130_fd_sc_hd__and2_1
Xclkbuf_4_9__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_9__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11802_ _11818_/B _11802_/B vssd1 vssd1 vccd1 vccd1 _11802_/X sky130_fd_sc_hd__and2_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15570_/A _15570_/B vssd1 vssd1 vccd1 vccd1 _15570_/X sky130_fd_sc_hd__xor2_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _17824_/Q _12781_/X _13944_/B vssd1 vssd1 vccd1 vccd1 _12782_/X sky130_fd_sc_hd__mux2_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _17723_/A0 _18371_/Q _14521_/S vssd1 vssd1 vccd1 vccd1 _18371_/D sky130_fd_sc_hd__mux2_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _18564_/Q _11741_/A2 _11769_/B1 _11732_/Y vssd1 vssd1 vccd1 vccd1 _11733_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _17238_/Y _17239_/X _17330_/A vssd1 vssd1 vccd1 vccd1 _19430_/D sky130_fd_sc_hd__a21oi_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14452_ _18592_/Q _14452_/B vssd1 vssd1 vccd1 vccd1 _18305_/D sky130_fd_sc_hd__and2_1
XFILLER_42_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11666_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11664_/X sky130_fd_sc_hd__and2_4
X_13403_ _12755_/A _12448_/C _13401_/Y _13402_/X _12762_/B vssd1 vssd1 vccd1 vccd1
+ _13403_/X sky130_fd_sc_hd__a221o_4
X_10615_ _10866_/S _10613_/X _10614_/X vssd1 vssd1 vccd1 vccd1 _10615_/X sky130_fd_sc_hd__o21a_1
X_17171_ _17285_/A _17171_/B vssd1 vssd1 vccd1 vccd1 _19408_/D sky130_fd_sc_hd__nor2_1
X_14383_ _18235_/Q _16557_/A0 _14383_/S vssd1 vssd1 vccd1 vccd1 _18235_/D sky130_fd_sc_hd__mux2_1
XFILLER_259_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11595_ _18874_/Q _18906_/Q _11598_/S vssd1 vssd1 vccd1 vccd1 _11595_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16122_ _16140_/A1 _16121_/Y _16142_/B1 vssd1 vssd1 vccd1 vccd1 _18763_/D sky130_fd_sc_hd__a21oi_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_259_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13334_ _17836_/Q _13844_/A2 _13844_/B1 _17868_/Q vssd1 vssd1 vccd1 vccd1 _13334_/X
+ sky130_fd_sc_hd__a22o_1
X_10546_ _10866_/S _18803_/Q _10613_/S vssd1 vssd1 vccd1 vccd1 _10546_/X sky130_fd_sc_hd__and3_1
XFILLER_143_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16053_ _18738_/Q _16069_/B _15854_/B vssd1 vssd1 vccd1 vccd1 _16053_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _13315_/S _13001_/Y _13264_/X vssd1 vssd1 vccd1 vccd1 _13265_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10477_ _10475_/X _10476_/X _10632_/S vssd1 vssd1 vccd1 vccd1 _10477_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15004_ _15002_/X _15003_/X _14714_/B vssd1 vssd1 vccd1 vccd1 _15004_/X sky130_fd_sc_hd__a21o_1
X_12216_ _17869_/Q _17870_/Q _12216_/C vssd1 vssd1 vccd1 vccd1 _12218_/B sky130_fd_sc_hd__and3_1
X_13196_ _14156_/A0 _13195_/X _09318_/B vssd1 vssd1 vccd1 vccd1 _13196_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_151_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ _17159_/A _12152_/C vssd1 vssd1 vccd1 vccd1 _12147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16955_ _19323_/Q _17202_/B _16963_/S vssd1 vssd1 vccd1 vccd1 _16956_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12078_ _17914_/Q _12086_/A2 _12077_/X _17419_/C1 vssd1 vssd1 vccd1 vccd1 _17816_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_256_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15906_ _18677_/Q _15906_/A2 _15906_/B1 _15905_/X vssd1 vssd1 vccd1 vccd1 _15906_/X
+ sky130_fd_sc_hd__a211o_1
X_11029_ _11512_/A1 _19636_/Q _18925_/Q _11513_/B2 vssd1 vssd1 vccd1 vccd1 _11029_/X
+ sky130_fd_sc_hd__a22o_1
X_16886_ _16898_/A1 _17930_/Q _16885_/X vssd1 vssd1 vccd1 vccd1 _17579_/A sky130_fd_sc_hd__o21a_4
XFILLER_265_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15837_ _15843_/A _15837_/B vssd1 vssd1 vccd1 vccd1 _15837_/Y sky130_fd_sc_hd__nand2_1
X_18625_ _19639_/CLK _18625_/D vssd1 vssd1 vccd1 vccd1 _18625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_252_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15768_ _15722_/B _15744_/B _15787_/A vssd1 vssd1 vccd1 vccd1 _15768_/Y sky130_fd_sc_hd__o21ai_1
X_18556_ _19638_/CLK _18556_/D vssd1 vssd1 vccd1 vccd1 _18556_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14719_ _14875_/B1 _14716_/X _14718_/Y _14928_/B1 vssd1 vssd1 vccd1 vccd1 _14720_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_17507_ _18124_/Q _17539_/C1 _17505_/X _17506_/X vssd1 vssd1 vccd1 vccd1 _17507_/X
+ sky130_fd_sc_hd__a22o_2
X_18487_ _19291_/CLK _18487_/D vssd1 vssd1 vccd1 vccd1 _18487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15699_ _18588_/Q _15800_/A2 _15691_/X _15698_/X _15718_/C1 vssd1 vssd1 vccd1 vccd1
+ _18588_/D sky130_fd_sc_hd__o221a_1
XFILLER_268_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_490 _18115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17438_ _17438_/A _17547_/B vssd1 vssd1 vccd1 vccd1 _17438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_15 _14879_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_26 _17172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_37 _09099_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 _12613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ _19482_/Q _17199_/B _17379_/S vssd1 vssd1 vccd1 vccd1 _17370_/B sky130_fd_sc_hd__mux2_1
XFILLER_158_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_59 _09995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19108_ _19140_/CLK _19108_/D vssd1 vssd1 vccd1 vccd1 _19108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19039_ _19138_/CLK _19039_/D vssd1 vssd1 vccd1 vccd1 _19039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_68_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19599_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_130_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09625_ _18848_/Q _18880_/Q _10313_/S vssd1 vssd1 vccd1 vccd1 _09625_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ _09611_/A _09555_/X _11790_/B vssd1 vssd1 vccd1 vccd1 _09556_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_271_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09487_ _09908_/A1 _09236_/A _09486_/X _09656_/B1 _18395_/Q vssd1 vssd1 vccd1 vccd1
+ _09487_/X sky130_fd_sc_hd__o32a_2
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10400_ _18558_/Q _18433_/Q _18042_/Q _18010_/Q _11462_/S _09136_/S vssd1 vssd1 vccd1
+ vccd1 _10400_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11380_ _10403_/S _11379_/X _11378_/X _09135_/S vssd1 vssd1 vccd1 vccd1 _11380_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_165_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10331_ _10336_/A _10330_/X _11466_/B1 vssd1 vssd1 vccd1 vccd1 _10331_/X sky130_fd_sc_hd__o21a_1
XFILLER_194_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10262_ _10262_/A1 _18232_/Q _09937_/S _18967_/Q vssd1 vssd1 vccd1 vccd1 _10262_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13050_ _13036_/X _13049_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _13051_/C sky130_fd_sc_hd__a21oi_1
XFILLER_152_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12001_ _17768_/Q _16470_/A0 _12021_/S vssd1 vssd1 vccd1 vccd1 _17768_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10193_ _10190_/X _10192_/X _10186_/X vssd1 vssd1 vccd1 vccd1 _10193_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_121_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1303 _16893_/A2 vssd1 vssd1 vccd1 vccd1 _16961_/A2 sky130_fd_sc_hd__buf_2
XFILLER_267_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1314 _11724_/Y vssd1 vssd1 vccd1 vccd1 _11759_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout1325 _09098_/Y vssd1 vssd1 vccd1 vccd1 _11237_/B1 sky130_fd_sc_hd__buf_4
Xfanout1336 _11459_/A1 vssd1 vssd1 vccd1 vccd1 _10336_/A sky130_fd_sc_hd__buf_4
XFILLER_238_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1347 _09463_/S vssd1 vssd1 vccd1 vccd1 _11161_/S sky130_fd_sc_hd__buf_8
XFILLER_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1358 _11224_/B vssd1 vssd1 vccd1 vccd1 _10838_/B sky130_fd_sc_hd__buf_4
XFILLER_120_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1369 _10929_/S vssd1 vssd1 vccd1 vccd1 _11302_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16740_ _16740_/A _16742_/B vssd1 vssd1 vccd1 vccd1 _16740_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13952_ _19327_/Q _13952_/A2 _13952_/B1 _13945_/X _13951_/X vssd1 vssd1 vccd1 vccd1
+ _13952_/Y sky130_fd_sc_hd__a2111oi_2
XFILLER_143_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12903_ _12448_/D _12899_/X _12902_/X _12871_/X vssd1 vssd1 vccd1 vccd1 _12903_/X
+ sky130_fd_sc_hd__a31o_1
X_16671_ _16776_/A _16673_/B vssd1 vssd1 vccd1 vccd1 _16671_/Y sky130_fd_sc_hd__nor2_1
XFILLER_262_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13883_ _19357_/Q _13883_/A2 _13883_/B1 _19485_/Q _13883_/C1 vssd1 vssd1 vccd1 vccd1
+ _13883_/X sky130_fd_sc_hd__a221o_1
XFILLER_234_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15622_ _18584_/Q _15621_/C _18585_/Q vssd1 vssd1 vccd1 vccd1 _15623_/C sky130_fd_sc_hd__a21oi_1
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18410_ _19148_/CLK _18410_/D vssd1 vssd1 vccd1 vccd1 _18410_/Q sky130_fd_sc_hd__dfxtp_1
X_19390_ _19458_/CLK _19390_/D vssd1 vssd1 vccd1 vccd1 _19390_/Q sky130_fd_sc_hd__dfxtp_2
X_12834_ _13315_/S _12833_/Y _13413_/B1 vssd1 vssd1 vccd1 vccd1 _12835_/B sky130_fd_sc_hd__a21o_1
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _19626_/CLK _18341_/D vssd1 vssd1 vccd1 vccd1 _18341_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15702_/A _15553_/B vssd1 vssd1 vccd1 vccd1 _15638_/A sky130_fd_sc_hd__xnor2_4
XFILLER_261_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _13257_/A _12765_/B vssd1 vssd1 vccd1 vccd1 _17920_/D sky130_fd_sc_hd__and2_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14504_ _16606_/A0 _18354_/Q _14516_/S vssd1 vssd1 vccd1 vccd1 _18354_/D sky130_fd_sc_hd__mux2_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18272_ _18272_/CLK _18272_/D vssd1 vssd1 vccd1 vccd1 _18272_/Q sky130_fd_sc_hd__dfxtp_2
X_11716_ _18531_/Q _18530_/Q vssd1 vssd1 vccd1 vccd1 _15835_/A sky130_fd_sc_hd__and2b_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15484_/A _15484_/B _15484_/C vssd1 vssd1 vccd1 vccd1 _15508_/B sky130_fd_sc_hd__nand3_2
XFILLER_30_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12696_ _12609_/B _12653_/B _13911_/A vssd1 vssd1 vccd1 vccd1 _12696_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17223_ _19425_/Q _17241_/B vssd1 vssd1 vccd1 vccd1 _17223_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14435_ _18574_/Q _17360_/A vssd1 vssd1 vccd1 vccd1 _18287_/D sky130_fd_sc_hd__and2_2
X_11647_ _11647_/A _11816_/A vssd1 vssd1 vccd1 vccd1 _11647_/X sky130_fd_sc_hd__or2_2
XFILLER_238_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 core_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17154_ _17157_/A _17581_/A vssd1 vssd1 vccd1 vccd1 _17448_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput24 core_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput35 core_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_2
X_14366_ _18218_/Q _16540_/A0 _14383_/S vssd1 vssd1 vccd1 vccd1 _18218_/D sky130_fd_sc_hd__mux2_1
X_11578_ _11574_/X _11577_/X _11578_/S vssd1 vssd1 vccd1 vccd1 _11579_/B sky130_fd_sc_hd__mux2_1
Xinput46 dout0[12] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_2
Xinput57 dout0[22] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_2
X_16105_ _18755_/Q _16137_/B vssd1 vssd1 vccd1 vccd1 _16105_/Y sky130_fd_sc_hd__nand2_1
Xinput68 dout0[32] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_2
X_13317_ _13316_/A _14155_/B _13316_/Y _13358_/A1 vssd1 vssd1 vccd1 vccd1 _13317_/X
+ sky130_fd_sc_hd__o211a_1
X_10529_ _17976_/Q _11295_/A2 _11216_/B1 vssd1 vssd1 vccd1 vccd1 _10529_/X sky130_fd_sc_hd__a21o_1
Xinput79 dout0[42] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_2
X_17085_ _19376_/Q _17115_/B vssd1 vssd1 vccd1 vccd1 _17085_/X sky130_fd_sc_hd__or2_1
XFILLER_128_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14297_ _17715_/A0 _18156_/Q _14305_/S vssd1 vssd1 vccd1 vccd1 _18156_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16036_ _15845_/A _16038_/A _18732_/Q vssd1 vssd1 vccd1 vccd1 _16036_/Y sky130_fd_sc_hd__o21ai_1
X_13248_ _15887_/A _12506_/X _13240_/X _13247_/X _12510_/X vssd1 vssd1 vccd1 vccd1
+ _13248_/X sky130_fd_sc_hd__o221a_1
XFILLER_170_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13179_ _13945_/B2 _13164_/X _13178_/X vssd1 vssd1 vccd1 vccd1 _13990_/B sky130_fd_sc_hd__a21oi_4
XFILLER_285_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17987_ _19148_/CLK _17987_/D vssd1 vssd1 vccd1 vccd1 _17987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1870 _08859_/Y vssd1 vssd1 vccd1 vccd1 fanout1870/X sky130_fd_sc_hd__buf_12
XFILLER_84_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16938_ _12482_/S _17943_/Q _16937_/X vssd1 vssd1 vccd1 vccd1 _17190_/B sky130_fd_sc_hd__o21a_4
XFILLER_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1881 fanout1905/X vssd1 vssd1 vccd1 vccd1 _17330_/A sky130_fd_sc_hd__buf_6
XFILLER_284_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1892 _16811_/A vssd1 vssd1 vccd1 vccd1 _12203_/A sky130_fd_sc_hd__buf_4
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16869_ _16848_/S _17926_/Q _16868_/X vssd1 vssd1 vccd1 vccd1 _17571_/A sky130_fd_sc_hd__o21a_4
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09410_ _10300_/S _09409_/X _11495_/B1 vssd1 vssd1 vccd1 vccd1 _09410_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18608_ _19216_/CLK _18608_/D vssd1 vssd1 vccd1 vccd1 _18608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19588_ _19588_/CLK _19588_/D vssd1 vssd1 vccd1 vccd1 _19588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09341_ _19203_/Q _19171_/Q _10099_/S vssd1 vssd1 vccd1 vccd1 _09341_/X sky130_fd_sc_hd__mux2_1
XFILLER_252_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18539_ _19591_/CLK _18539_/D vssd1 vssd1 vccd1 vccd1 _18539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_186_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19092_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_279_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09272_ _09272_/A1 _19140_/Q _09252_/S _19108_/Q _10408_/S vssd1 vssd1 vccd1 vccd1
+ _09272_/X sky130_fd_sc_hd__o221a_1
XFILLER_179_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_115_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19286_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ _18268_/Q _18200_/Q vssd1 vssd1 vccd1 vccd1 _08987_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09608_ _09608_/A _09608_/B vssd1 vssd1 vccd1 vccd1 _09608_/Y sky130_fd_sc_hd__nand2_2
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10880_ _11355_/A1 _10879_/X _11286_/B1 vssd1 vssd1 vccd1 vccd1 _10880_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ _18849_/Q _18881_/Q _09539_/S vssd1 vssd1 vccd1 vccd1 _09539_/X sky130_fd_sc_hd__mux2_1
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12550_ _13945_/B2 _12498_/X _12549_/X vssd1 vssd1 vccd1 vccd1 _12550_/X sky130_fd_sc_hd__a21o_4
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11501_ _09967_/S _11500_/X _11501_/B1 vssd1 vssd1 vccd1 vccd1 _11501_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ _12501_/A _12501_/B _12502_/A vssd1 vssd1 vccd1 vccd1 _12491_/A sky130_fd_sc_hd__or3_1
XFILLER_169_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14220_ _14220_/A _14224_/B vssd1 vssd1 vccd1 vccd1 _14220_/Y sky130_fd_sc_hd__nand2_1
X_11432_ _18249_/Q _18824_/Q _18452_/Q _18353_/Q _11513_/B2 _11510_/S1 vssd1 vssd1
+ vccd1 vccd1 _11433_/B sky130_fd_sc_hd__mux4_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _14151_/A _14151_/B _14151_/C _14151_/D vssd1 vssd1 vccd1 vccd1 _14153_/C
+ sky130_fd_sc_hd__nor4_4
X_11363_ _11358_/Y _11362_/Y _11621_/C1 vssd1 vssd1 vccd1 vccd1 _11363_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13102_ _17830_/Q _13164_/A2 _13164_/B1 _17862_/Q vssd1 vssd1 vccd1 vccd1 _13102_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10314_ _18466_/Q _18367_/Q _10687_/S vssd1 vssd1 vccd1 vccd1 _10314_/X sky130_fd_sc_hd__mux2_1
X_14082_ _16532_/A0 _18022_/Q _14104_/S vssd1 vssd1 vccd1 vccd1 _18022_/D sky130_fd_sc_hd__mux2_1
X_11294_ _12626_/A vssd1 vssd1 vccd1 vccd1 _13411_/A sky130_fd_sc_hd__inv_4
XFILLER_279_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17910_ _19140_/CLK _17910_/D vssd1 vssd1 vccd1 vccd1 _17910_/Q sky130_fd_sc_hd__dfxtp_1
X_13033_ _13033_/A _13033_/B vssd1 vssd1 vccd1 vccd1 _13083_/C sky130_fd_sc_hd__nand2_1
XFILLER_112_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10245_ _19063_/Q _19031_/Q _10253_/C vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18890_ _19601_/CLK _18890_/D vssd1 vssd1 vccd1 vccd1 _18890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_279_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1100 _08882_/Y vssd1 vssd1 vccd1 vccd1 _17546_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_133_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1111 _12455_/Y vssd1 vssd1 vccd1 vccd1 _13929_/A1 sky130_fd_sc_hd__buf_6
X_10176_ _18872_/Q _18904_/Q _10176_/S vssd1 vssd1 vccd1 vccd1 _10176_/X sky130_fd_sc_hd__mux2_1
X_17841_ _19363_/CLK _17841_/D vssd1 vssd1 vccd1 vccd1 _17841_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1122 _13791_/A vssd1 vssd1 vccd1 vccd1 _13462_/A sky130_fd_sc_hd__buf_6
XFILLER_267_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1133 _13936_/B2 vssd1 vssd1 vccd1 vccd1 _12761_/B sky130_fd_sc_hd__buf_4
Xfanout1144 _10239_/A vssd1 vssd1 vccd1 vccd1 _11452_/A sky130_fd_sc_hd__buf_8
XFILLER_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1155 _16002_/C1 vssd1 vssd1 vccd1 vccd1 _15976_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1166 _15852_/X vssd1 vssd1 vccd1 vccd1 _15948_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_254_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14984_ _14982_/X _14983_/X _14995_/A1 vssd1 vssd1 vccd1 vccd1 _14984_/X sky130_fd_sc_hd__a21o_1
X_17772_ _19600_/CLK _17772_/D vssd1 vssd1 vccd1 vccd1 _17772_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1177 _13260_/Y vssd1 vssd1 vccd1 vccd1 _13892_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1188 _08948_/B vssd1 vssd1 vccd1 vccd1 _11451_/A2 sky130_fd_sc_hd__buf_6
XFILLER_248_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1199 _12837_/X vssd1 vssd1 vccd1 vccd1 _13797_/A0 sky130_fd_sc_hd__buf_6
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19511_ _19531_/CLK _19511_/D vssd1 vssd1 vccd1 vccd1 _19511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16723_ _19260_/Q _19259_/Q _16723_/C vssd1 vssd1 vccd1 vccd1 _16729_/C sky130_fd_sc_hd__and3_1
X_13935_ _13969_/B _13935_/B vssd1 vssd1 vccd1 vccd1 _13935_/Y sky130_fd_sc_hd__nand2_2
XFILLER_35_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16654_ _19240_/Q _16658_/C vssd1 vssd1 vccd1 vccd1 _16661_/C sky130_fd_sc_hd__and2_1
X_19442_ _19519_/CLK _19442_/D vssd1 vssd1 vccd1 vccd1 _19442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_262_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13866_ _13289_/A _13857_/X _13858_/Y _17531_/A _13294_/A vssd1 vssd1 vccd1 vccd1
+ _13866_/X sky130_fd_sc_hd__o32a_1
XFILLER_250_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15605_ _15690_/A _15603_/Y _15604_/X _15751_/A vssd1 vssd1 vccd1 vccd1 _15605_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_262_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12817_ _12817_/A vssd1 vssd1 vccd1 vccd1 _12817_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19373_ _19470_/CLK _19373_/D vssd1 vssd1 vccd1 vccd1 _19373_/Q sky130_fd_sc_hd__dfxtp_1
X_16585_ _16618_/A0 _19189_/Q _16585_/S vssd1 vssd1 vccd1 vccd1 _19189_/D sky130_fd_sc_hd__mux2_1
X_13797_ _13797_/A0 _12756_/Y _13797_/S vssd1 vssd1 vccd1 vccd1 _13797_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15536_ _15554_/B _15536_/B vssd1 vssd1 vccd1 vccd1 _15536_/Y sky130_fd_sc_hd__xnor2_1
X_18324_ _18613_/CLK _18324_/D vssd1 vssd1 vccd1 vccd1 _18324_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12748_/A vssd1 vssd1 vccd1 vccd1 _12748_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18255_ _19573_/CLK _18255_/D vssd1 vssd1 vccd1 vccd1 _18255_/Q sky130_fd_sc_hd__dfxtp_1
X_15467_ _15512_/C _15467_/B vssd1 vssd1 vccd1 vccd1 _15467_/X sky130_fd_sc_hd__or2_1
X_12679_ _10982_/Y _12625_/B _12704_/S vssd1 vssd1 vccd1 vccd1 _12680_/A sky130_fd_sc_hd__mux2_4
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17206_ _19420_/Q fanout533/X _17205_/Y _17119_/B vssd1 vssd1 vccd1 vccd1 _17207_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14418_ _19227_/Q _15014_/B _18274_/D vssd1 vssd1 vccd1 vccd1 _18269_/D sky130_fd_sc_hd__and3_1
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18186_ _19639_/CLK _18186_/D vssd1 vssd1 vccd1 vccd1 _18186_/Q sky130_fd_sc_hd__dfxtp_1
X_15398_ _15398_/A _15398_/B vssd1 vssd1 vccd1 vccd1 _15399_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17137_ _19397_/Q fanout534/X _17418_/A _17212_/B2 vssd1 vssd1 vccd1 vccd1 _17138_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14349_ _14430_/B _14349_/B vssd1 vssd1 vccd1 vccd1 _18203_/D sky130_fd_sc_hd__and2_2
XFILLER_7_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17068_ _17573_/A _17114_/A2 _17067_/X _17559_/A vssd1 vssd1 vccd1 vccd1 _19367_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16019_ _18725_/Q _16019_/A2 _16018_/X _14197_/A vssd1 vssd1 vccd1 vccd1 _18725_/D
+ sky130_fd_sc_hd__o211a_1
X_08910_ _08940_/B _08929_/B vssd1 vssd1 vccd1 vccd1 _08939_/A sky130_fd_sc_hd__nor2_8
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _11189_/A _09882_/X _09881_/X _11198_/S vssd1 vssd1 vccd1 vccd1 _09890_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_258_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _17914_/Q vssd1 vssd1 vccd1 vccd1 _08841_/Y sky130_fd_sc_hd__inv_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09324_ _09012_/A _09236_/A _09323_/X _09656_/B1 _18389_/Q vssd1 vssd1 vccd1 vccd1
+ _09325_/D sky130_fd_sc_hd__o32a_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09255_ _19204_/Q _19172_/Q _11395_/C vssd1 vssd1 vccd1 vccd1 _09255_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09186_ _09186_/A _09186_/B vssd1 vssd1 vccd1 vccd1 _09186_/X sky130_fd_sc_hd__and2_1
XFILLER_194_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_83_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18881_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_175_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19025_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10030_ _11284_/A1 _19195_/Q _19163_/Q _11617_/S _10030_/C1 vssd1 vssd1 vccd1 vccd1
+ _10030_/X sky130_fd_sc_hd__a221o_1
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput203 localMemory_wb_adr_i[21] vssd1 vssd1 vccd1 vccd1 _12269_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput214 localMemory_wb_cyc_i vssd1 vssd1 vccd1 vccd1 _15013_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_102_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput225 localMemory_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input225/X sky130_fd_sc_hd__clkbuf_16
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput236 localMemory_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 input236/X sky130_fd_sc_hd__clkbuf_16
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput247 localMemory_wb_sel_i[0] vssd1 vssd1 vccd1 vccd1 input247/X sky130_fd_sc_hd__clkbuf_2
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput258 manufacturerID[4] vssd1 vssd1 vccd1 vccd1 _15869_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput269 partID[14] vssd1 vssd1 vccd1 vccd1 input269/X sky130_fd_sc_hd__clkbuf_2
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ _18741_/Q _11981_/B vssd1 vssd1 vccd1 vccd1 _16069_/B sky130_fd_sc_hd__or2_2
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13720_ _19352_/Q _13883_/A2 _13883_/B1 _19480_/Q _13883_/C1 vssd1 vssd1 vccd1 vccd1
+ _13720_/X sky130_fd_sc_hd__a221o_1
X_10932_ _11327_/S _19182_/Q _10940_/S vssd1 vssd1 vccd1 vccd1 _10932_/X sky130_fd_sc_hd__and3_1
XFILLER_244_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13651_ _17877_/Q _13747_/A2 _13650_/X _13682_/B2 vssd1 vssd1 vccd1 vccd1 _13651_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_271_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10863_ _11577_/S _10862_/X _11328_/S vssd1 vssd1 vccd1 vccd1 _10863_/X sky130_fd_sc_hd__a21o_1
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12602_ _12602_/A _12602_/B vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__or2_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _16470_/A0 _18981_/Q _16390_/S vssd1 vssd1 vccd1 vccd1 _18981_/D sky130_fd_sc_hd__mux2_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _17843_/Q _13744_/A2 _13744_/B1 _17875_/Q vssd1 vssd1 vccd1 vccd1 _13582_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10794_ _10471_/S _11135_/S _11181_/B1 _10793_/Y vssd1 vssd1 vccd1 vccd1 _10832_/A
+ sky130_fd_sc_hd__o22a_2
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15319_/Y _15321_/B vssd1 vssd1 vccd1 vccd1 _15324_/A sky130_fd_sc_hd__nand2b_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12533_ _13165_/B _12584_/A vssd1 vssd1 vccd1 vccd1 _12533_/Y sky130_fd_sc_hd__nor2_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18040_ _19638_/CLK _18040_/D vssd1 vssd1 vccd1 vccd1 _18040_/Q sky130_fd_sc_hd__dfxtp_1
X_15252_ _19463_/Q _19397_/Q vssd1 vssd1 vccd1 vccd1 _15254_/A sky130_fd_sc_hd__xnor2_1
XFILLER_200_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12464_ _12482_/S _14680_/B vssd1 vssd1 vccd1 vccd1 _16839_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14203_ _14203_/A _14203_/B vssd1 vssd1 vccd1 vccd1 _18099_/D sky130_fd_sc_hd__and2_1
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11415_ _11512_/A1 _18320_/Q _17771_/Q _11426_/B2 vssd1 vssd1 vccd1 vccd1 _11415_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15183_ _15224_/C _15183_/B vssd1 vssd1 vccd1 vccd1 _15183_/X sky130_fd_sc_hd__or2_1
X_12395_ _17906_/Q _12408_/B _12394_/Y _13981_/C1 vssd1 vssd1 vccd1 vccd1 _17906_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14134_ _17684_/A0 _18073_/Q _14140_/S vssd1 vssd1 vccd1 vccd1 _18073_/D sky130_fd_sc_hd__mux2_1
X_11346_ _11344_/X _11345_/X _11361_/S vssd1 vssd1 vccd1 vccd1 _11346_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14065_ _17682_/A0 _18007_/Q _14073_/S vssd1 vssd1 vccd1 vccd1 _18007_/D sky130_fd_sc_hd__mux2_1
X_18942_ _19134_/CLK _18942_/D vssd1 vssd1 vccd1 vccd1 _18942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11277_ _11277_/A1 _19114_/Q _19146_/Q _11617_/S vssd1 vssd1 vccd1 vccd1 _11277_/X
+ sky130_fd_sc_hd__a22o_1
X_13016_ _19397_/Q _12570_/A _13244_/B1 vssd1 vssd1 vccd1 vccd1 _13016_/X sky130_fd_sc_hd__a21o_1
X_10228_ _11417_/B1 _10210_/X _10211_/X _10221_/X _10227_/X vssd1 vssd1 vccd1 vccd1
+ _10228_/X sky130_fd_sc_hd__o32a_4
X_18873_ _19193_/CLK _18873_/D vssd1 vssd1 vccd1 vccd1 _18873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17824_ _18761_/CLK _17824_/D vssd1 vssd1 vccd1 vccd1 _17824_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10159_ _10159_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _13913_/A sky130_fd_sc_hd__nor2_1
XFILLER_95_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17755_ _18655_/Q vssd1 vssd1 vccd1 vccd1 _18655_/D sky130_fd_sc_hd__clkbuf_2
X_14967_ input62/X input97/X _15007_/S vssd1 vssd1 vccd1 vccd1 _14968_/A sky130_fd_sc_hd__mux2_2
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16706_ _19255_/Q _16706_/B vssd1 vssd1 vccd1 vccd1 _16713_/C sky130_fd_sc_hd__and2_1
X_13918_ _17853_/Q _13942_/A2 _13942_/B1 _17885_/Q vssd1 vssd1 vccd1 vccd1 _13918_/X
+ sky130_fd_sc_hd__a22o_1
X_17686_ _17686_/A0 _19613_/Q _17689_/S vssd1 vssd1 vccd1 vccd1 _19613_/D sky130_fd_sc_hd__mux2_1
XFILLER_223_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14898_ _14979_/A1 _18271_/Q _14897_/Y _14918_/B1 vssd1 vssd1 vccd1 vccd1 _14898_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_251_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19425_ _19525_/CLK _19425_/D vssd1 vssd1 vccd1 vccd1 _19425_/Q sky130_fd_sc_hd__dfxtp_1
X_16637_ _19234_/Q _16677_/A _19235_/Q vssd1 vssd1 vccd1 vccd1 _16639_/B sky130_fd_sc_hd__a21oi_1
X_13849_ _19518_/Q _13947_/A2 _13947_/B1 _13848_/X vssd1 vssd1 vccd1 vccd1 _13849_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19356_ _19542_/CLK _19356_/D vssd1 vssd1 vccd1 vccd1 _19356_/Q sky130_fd_sc_hd__dfxtp_1
X_16568_ _17668_/A0 _19172_/Q _16589_/S vssd1 vssd1 vccd1 vccd1 _19172_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18307_ _19586_/CLK _18307_/D vssd1 vssd1 vccd1 vccd1 _18307_/Q sky130_fd_sc_hd__dfxtp_1
X_15519_ _19474_/Q _19408_/Q vssd1 vssd1 vccd1 vccd1 _15519_/Y sky130_fd_sc_hd__nor2_1
X_19287_ _19291_/CLK _19287_/D vssd1 vssd1 vccd1 vccd1 _19287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16499_ _16532_/A0 _19105_/Q _16515_/S vssd1 vssd1 vccd1 vccd1 _19105_/D sky130_fd_sc_hd__mux2_1
XFILLER_198_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09040_ _09043_/A _09032_/B _08913_/X _08939_/A vssd1 vssd1 vccd1 vccd1 _09042_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_191_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18238_ _19133_/CLK _18238_/D vssd1 vssd1 vccd1 vccd1 _18238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18169_ _19138_/CLK _18169_/D vssd1 vssd1 vccd1 vccd1 _18169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09942_ _10194_/C1 _09980_/A2 _09941_/X _11023_/B1 vssd1 vssd1 vccd1 vccd1 _11785_/B
+ sky130_fd_sc_hd__o211ai_4
Xfanout904 _16458_/S vssd1 vssd1 vccd1 vccd1 _16453_/S sky130_fd_sc_hd__buf_12
XFILLER_132_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout915 _16359_/X vssd1 vssd1 vccd1 vccd1 _16388_/S sky130_fd_sc_hd__buf_8
Xfanout926 _16212_/S vssd1 vssd1 vccd1 vccd1 _16222_/S sky130_fd_sc_hd__buf_12
XFILLER_86_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout937 _14982_/B vssd1 vssd1 vccd1 vccd1 _14911_/B sky130_fd_sc_hd__clkbuf_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _09873_/A1 _19620_/Q _18909_/Q _10054_/S _15481_/A vssd1 vssd1 vccd1 vccd1
+ _09873_/X sky130_fd_sc_hd__a221o_1
Xfanout948 _14670_/Y vssd1 vssd1 vccd1 vccd1 _14995_/A1 sky130_fd_sc_hd__buf_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout959 _14521_/S vssd1 vssd1 vccd1 vccd1 _14517_/S sky130_fd_sc_hd__buf_12
XFILLER_140_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _18774_/Q vssd1 vssd1 vccd1 vccd1 _16143_/C sky130_fd_sc_hd__inv_2
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 _18113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_130_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19502_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_319 _18104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09307_ _11498_/A1 _18213_/Q _09306_/S _18948_/Q _09374_/S vssd1 vssd1 vccd1 vccd1
+ _09307_/X sky130_fd_sc_hd__o221a_1
XFILLER_167_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09238_ _09901_/A vssd1 vssd1 vccd1 vccd1 _09238_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09169_ _09167_/X _09168_/X _10169_/S vssd1 vssd1 vccd1 vccd1 _09169_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _09718_/S _11199_/X _08903_/A vssd1 vssd1 vccd1 vccd1 _11200_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12180_ _17856_/Q _12178_/B _12179_/Y vssd1 vssd1 vccd1 vccd1 _17856_/D sky130_fd_sc_hd__o21a_1
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11131_ _11131_/A _11131_/B _11131_/C vssd1 vssd1 vccd1 vccd1 _11131_/X sky130_fd_sc_hd__or3_1
XFILLER_268_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ _13535_/S _11062_/B vssd1 vssd1 vccd1 vccd1 _12593_/A sky130_fd_sc_hd__nor2_8
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10013_ _19618_/Q _18907_/Q _11581_/S vssd1 vssd1 vccd1 vccd1 _10013_/X sky130_fd_sc_hd__mux2_1
X_15870_ _18665_/Q _15853_/Y _15903_/B1 vssd1 vssd1 vccd1 vccd1 _15870_/X sky130_fd_sc_hd__a21o_1
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _18114_/Q _14994_/B vssd1 vssd1 vccd1 vccd1 _14821_/X sky130_fd_sc_hd__or2_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _14750_/X _14751_/X _14964_/B1 vssd1 vssd1 vccd1 vccd1 _14752_/X sky130_fd_sc_hd__a21o_1
X_17540_ _18130_/Q _08883_/A _17540_/B1 _17539_/X vssd1 vssd1 vccd1 vccd1 _17540_/Y
+ sky130_fd_sc_hd__o211ai_2
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _18510_/Q _11720_/X _11914_/X _11968_/B2 vssd1 vssd1 vccd1 vccd1 _11964_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_245_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _13968_/A1 _13694_/X _13702_/X _13323_/B vssd1 vssd1 vccd1 vccd1 _13703_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17471_ _18578_/Q _17544_/A _08883_/A vssd1 vssd1 vccd1 vccd1 _17471_/X sky130_fd_sc_hd__o21a_1
X_10915_ _19086_/Q _11581_/S _10914_/X _11559_/S1 vssd1 vssd1 vccd1 vccd1 _10915_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_260_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14683_ _14683_/A _14683_/B vssd1 vssd1 vccd1 vccd1 _14683_/X sky130_fd_sc_hd__and2_2
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11895_ _10196_/B _11845_/B _11952_/A2 vssd1 vssd1 vccd1 vccd1 _11899_/B sky130_fd_sc_hd__o21ai_2
XFILLER_233_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19210_ _19640_/CLK _19210_/D vssd1 vssd1 vccd1 vccd1 _19210_/Q sky130_fd_sc_hd__dfxtp_1
X_16422_ _16455_/A1 _19031_/Q _16424_/S vssd1 vssd1 vccd1 vccd1 _19031_/D sky130_fd_sc_hd__mux2_1
X_13634_ _19317_/Q _13174_/A _13722_/B1 _13627_/X _13633_/X vssd1 vssd1 vccd1 vccd1
+ _13634_/Y sky130_fd_sc_hd__a2111oi_2
XFILLER_220_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10846_ _18427_/Q _11300_/B _10845_/X _10557_/S vssd1 vssd1 vccd1 vccd1 _10846_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16353_ _18965_/Q _17685_/A0 _16357_/S vssd1 vssd1 vccd1 vccd1 _18965_/D sky130_fd_sc_hd__mux2_1
X_19141_ _19604_/CLK _19141_/D vssd1 vssd1 vccd1 vccd1 _19141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13565_ _13622_/A _13566_/A _13564_/X vssd1 vssd1 vccd1 vccd1 _13565_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10777_ _11572_/A1 _19575_/Q _10853_/S _19607_/Q vssd1 vssd1 vccd1 vccd1 _10777_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15304_ _15304_/A1 _13236_/Y _15381_/A3 _15303_/X vssd1 vssd1 vccd1 vccd1 _15304_/X
+ sky130_fd_sc_hd__a31o_1
X_12516_ _12768_/A _12584_/A vssd1 vssd1 vccd1 vccd1 _12516_/Y sky130_fd_sc_hd__nor2_1
X_19072_ _19211_/CLK _19072_/D vssd1 vssd1 vccd1 vccd1 _19072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16284_ _17715_/A0 _18898_/Q _16292_/S vssd1 vssd1 vccd1 vccd1 _18898_/D sky130_fd_sc_hd__mux2_1
X_13496_ _17872_/Q _13747_/A2 _13495_/X _13747_/B2 vssd1 vssd1 vccd1 vccd1 _13496_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18023_ _18880_/CLK _18023_/D vssd1 vssd1 vccd1 vccd1 _18023_/Q sky130_fd_sc_hd__dfxtp_1
X_15235_ _17389_/B1 _15234_/X _15424_/C1 vssd1 vssd1 vccd1 vccd1 _15235_/X sky130_fd_sc_hd__a21o_1
X_12447_ _12443_/D _12446_/X _12445_/A vssd1 vssd1 vccd1 vccd1 _12447_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_246_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15166_ _15166_/A _15166_/B vssd1 vssd1 vccd1 vccd1 _15167_/B sky130_fd_sc_hd__nor2_1
X_12378_ _18386_/Q _12429_/B1 _09567_/B _08858_/A vssd1 vssd1 vccd1 vccd1 _12379_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_153_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14117_ _16501_/A0 _18056_/Q _14139_/S vssd1 vssd1 vccd1 vccd1 _18056_/D sky130_fd_sc_hd__mux2_1
X_11329_ _11303_/X _11306_/X _10399_/A vssd1 vssd1 vccd1 vccd1 _11329_/X sky130_fd_sc_hd__a21o_1
X_15097_ _19378_/Q _15086_/B input179/X _15096_/X vssd1 vssd1 vccd1 vccd1 _15097_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18925_ _19636_/CLK _18925_/D vssd1 vssd1 vccd1 vccd1 _18925_/Q sky130_fd_sc_hd__dfxtp_1
X_14048_ _15808_/A1 _17990_/Q _14070_/S vssd1 vssd1 vccd1 vccd1 _17990_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18856_ _19208_/CLK _18856_/D vssd1 vssd1 vccd1 vccd1 _18856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17807_ _17814_/CLK _17807_/D vssd1 vssd1 vccd1 vccd1 _17807_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18787_ _19626_/CLK _18787_/D vssd1 vssd1 vccd1 vccd1 _18787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_283_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15999_ _18715_/Q _16005_/A2 _15998_/X _14205_/A vssd1 vssd1 vccd1 vccd1 _18715_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_282_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17738_ _18638_/Q vssd1 vssd1 vccd1 vccd1 _18638_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_36_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17669_ _17669_/A0 _19596_/Q _17689_/S vssd1 vssd1 vccd1 vccd1 _19596_/D sky130_fd_sc_hd__mux2_1
XFILLER_224_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19408_ _19540_/CLK _19408_/D vssd1 vssd1 vccd1 vccd1 _19408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19339_ _19534_/CLK _19339_/D vssd1 vssd1 vccd1 vccd1 _19339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09023_ _09043_/A _11218_/B _08990_/X vssd1 vssd1 vccd1 vccd1 _09023_/X sky130_fd_sc_hd__o21ba_1
XFILLER_176_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout701 _12544_/Y vssd1 vssd1 vccd1 vccd1 _13943_/A2 sky130_fd_sc_hd__buf_4
XFILLER_160_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout712 _12542_/Y vssd1 vssd1 vccd1 vccd1 _13115_/C1 sky130_fd_sc_hd__buf_4
X_09925_ _18237_/Q _18812_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _09925_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout723 _12497_/Y vssd1 vssd1 vccd1 vccd1 _13164_/B1 sky130_fd_sc_hd__buf_2
XFILLER_132_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout734 _11375_/X vssd1 vssd1 vccd1 vccd1 _16539_/A0 sky130_fd_sc_hd__buf_2
Xfanout745 _09947_/Y vssd1 vssd1 vccd1 vccd1 _12878_/S sky130_fd_sc_hd__buf_4
XFILLER_219_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout756 _09735_/A vssd1 vssd1 vccd1 vccd1 _12739_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout767 _17723_/S vssd1 vssd1 vccd1 vccd1 _17722_/S sky130_fd_sc_hd__clkbuf_16
X_09856_ _10707_/A _09851_/X _09855_/X _09534_/S vssd1 vssd1 vccd1 vccd1 _09856_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout778 _16619_/S vssd1 vssd1 vccd1 vccd1 _16622_/S sky130_fd_sc_hd__buf_12
XFILLER_213_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout789 _16492_/Y vssd1 vssd1 vccd1 vccd1 _16524_/S sky130_fd_sc_hd__buf_12
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_8__f_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_8__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _11284_/A1 _18136_/Q _18782_/Q _09797_/S _08899_/A vssd1 vssd1 vccd1 vccd1
+ _09787_/X sky130_fd_sc_hd__a221o_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_105 _11719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _11846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_127 _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _11836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _11868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10700_ _11250_/A1 _17780_/Q _11171_/S _18329_/Q vssd1 vssd1 vccd1 vccd1 _10700_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _13351_/A _11680_/B vssd1 vssd1 vccd1 vccd1 _13366_/B sky130_fd_sc_hd__xor2_4
XFILLER_241_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10631_ _10850_/A1 _19154_/Q _10634_/S0 _19122_/Q vssd1 vssd1 vccd1 vccd1 _10631_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13350_ _11681_/A _13311_/B _12625_/Y vssd1 vssd1 vccd1 vccd1 _13351_/B sky130_fd_sc_hd__a21oi_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10562_ _10623_/A _10540_/X _10548_/Y _10554_/Y _10561_/Y vssd1 vssd1 vccd1 vccd1
+ _10562_/X sky130_fd_sc_hd__a32o_1
XFILLER_195_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _14675_/C _12301_/B _14675_/B vssd1 vssd1 vccd1 vccd1 _12308_/B sky130_fd_sc_hd__or3b_1
XFILLER_10_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13281_ _19371_/Q _13280_/X _13925_/S vssd1 vssd1 vccd1 vccd1 _13281_/X sky130_fd_sc_hd__mux2_2
XFILLER_182_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10493_ _10491_/X _10492_/X _10643_/S vssd1 vssd1 vccd1 vccd1 _10493_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15020_ _18509_/Q input209/X _15024_/S vssd1 vssd1 vccd1 vccd1 _18509_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12232_ _17875_/Q _17876_/Q _12232_/C vssd1 vssd1 vccd1 vccd1 _12234_/B sky130_fd_sc_hd__and3_1
XFILLER_170_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12163_ _12243_/A _12168_/C vssd1 vssd1 vccd1 vccd1 _12163_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11114_ _11284_/A1 _19116_/Q _19148_/Q _09801_/S vssd1 vssd1 vccd1 vccd1 _11114_/X
+ sky130_fd_sc_hd__a22o_1
X_12094_ _17823_/Q _17824_/Q _17825_/Q vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__a21oi_1
X_16971_ _19327_/Q _17214_/B _16971_/S vssd1 vssd1 vccd1 vccd1 _16972_/B sky130_fd_sc_hd__mux2_1
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18710_ _18713_/CLK _18710_/D vssd1 vssd1 vccd1 vccd1 _18710_/Q sky130_fd_sc_hd__dfxtp_1
X_15922_ _18683_/Q _15943_/A2 _15921_/X _15946_/C1 vssd1 vssd1 vccd1 vccd1 _18683_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_277_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11045_ _09374_/S _11042_/X _11044_/X vssd1 vssd1 vccd1 vccd1 _11053_/B sky130_fd_sc_hd__a21oi_1
XFILLER_89_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18641_ _19586_/CLK _18641_/D vssd1 vssd1 vccd1 vccd1 _18641_/Q sky130_fd_sc_hd__dfxtp_4
X_15853_ _15853_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15853_/Y sky130_fd_sc_hd__nand2_4
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14804_ input45/X input80/X _14844_/S vssd1 vssd1 vccd1 vccd1 _14805_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18572_ _19465_/CLK _18572_/D vssd1 vssd1 vccd1 vccd1 _18572_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_218_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ _15767_/Y _15770_/B _15766_/A vssd1 vssd1 vccd1 vccd1 _15788_/A sky130_fd_sc_hd__o21ai_1
X_12996_ _12994_/A _12995_/X _13135_/S vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__mux2_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _19516_/Q _17523_/B vssd1 vssd1 vccd1 vccd1 _17523_/X sky130_fd_sc_hd__or2_1
XFILLER_217_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11947_ _14667_/A1 _11890_/B _11890_/C _11953_/A2 input234/X vssd1 vssd1 vccd1 vccd1
+ _11947_/X sky130_fd_sc_hd__a32o_4
X_14735_ _14214_/A _14801_/B _14690_/Y _14734_/X vssd1 vssd1 vccd1 vccd1 _14735_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14666_ _14667_/A1 _14417_/B _14665_/X vssd1 vssd1 vccd1 vccd1 _14666_/X sky130_fd_sc_hd__a21o_2
X_17454_ _19502_/Q _17453_/B _17452_/X _17453_/Y _17559_/A vssd1 vssd1 vccd1 vccd1
+ _19502_/D sky130_fd_sc_hd__o221a_1
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11878_ _11899_/A _11878_/B _11878_/C vssd1 vssd1 vccd1 vccd1 _11878_/X sky130_fd_sc_hd__and3_4
XFILLER_189_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16405_ _09105_/A _19014_/Q _16424_/S vssd1 vssd1 vccd1 vccd1 _19014_/D sky130_fd_sc_hd__mux2_1
X_13617_ _13761_/B _14149_/A _13892_/B1 vssd1 vssd1 vccd1 vccd1 _13617_/Y sky130_fd_sc_hd__a21oi_1
X_10829_ _18122_/Q _10828_/Y _10905_/S vssd1 vssd1 vccd1 vccd1 _12640_/B sky130_fd_sc_hd__mux2_4
XFILLER_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14597_ _08884_/X _09083_/A _11730_/Y _14594_/X vssd1 vssd1 vccd1 vccd1 _14597_/X
+ sky130_fd_sc_hd__o31a_1
X_17385_ _19489_/Q _12460_/A _15411_/B _17384_/X _14430_/B vssd1 vssd1 vccd1 vccd1
+ _19488_/D sky130_fd_sc_hd__o311a_1
X_19124_ _19620_/CLK _19124_/D vssd1 vssd1 vccd1 vccd1 _19124_/Q sky130_fd_sc_hd__dfxtp_1
X_16336_ _18948_/Q _16535_/A0 _16357_/S vssd1 vssd1 vccd1 vccd1 _18948_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13548_ _15526_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13548_/X sky130_fd_sc_hd__or2_2
XFILLER_173_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16267_ _17698_/A0 _18881_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _18881_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19055_ _19055_/CLK _19055_/D vssd1 vssd1 vccd1 vccd1 _19055_/Q sky130_fd_sc_hd__dfxtp_1
X_13479_ _18118_/Q _14238_/A _13479_/C vssd1 vssd1 vccd1 vccd1 _13541_/B sky130_fd_sc_hd__and3_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18006_ _19645_/CLK _18006_/D vssd1 vssd1 vccd1 vccd1 _18006_/Q sky130_fd_sc_hd__dfxtp_1
X_15218_ _12318_/A _15215_/Y _15216_/X _15369_/A _17914_/Q vssd1 vssd1 vccd1 vccd1
+ _15218_/Y sky130_fd_sc_hd__o2111ai_4
Xoutput304 _19653_/X vssd1 vssd1 vccd1 vccd1 clk1 sky130_fd_sc_hd__clkbuf_2
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16198_ _17695_/A0 _18814_/Q _16226_/S vssd1 vssd1 vccd1 vccd1 _18814_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput315 _11763_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[19] sky130_fd_sc_hd__buf_4
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput326 _11736_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[3] sky130_fd_sc_hd__buf_4
Xoutput337 _11822_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[12] sky130_fd_sc_hd__buf_4
X_15149_ _15135_/A _15135_/B _15138_/C vssd1 vssd1 vccd1 vccd1 _15149_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_236_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput348 _11868_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[22] sky130_fd_sc_hd__buf_4
Xoutput359 _11792_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[3] sky130_fd_sc_hd__buf_4
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09710_ _10742_/A1 _09704_/X _09705_/X vssd1 vssd1 vccd1 vccd1 _09710_/X sky130_fd_sc_hd__o21a_1
XFILLER_256_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18908_ _19619_/CLK _18908_/D vssd1 vssd1 vccd1 vccd1 _18908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09641_ _10180_/A _09635_/X _09640_/X _09617_/Y _09634_/Y vssd1 vssd1 vccd1 vccd1
+ _09641_/X sky130_fd_sc_hd__a32o_4
XFILLER_283_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18839_ _19646_/CLK _18839_/D vssd1 vssd1 vccd1 vccd1 _18839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09572_ _09908_/A1 _09236_/A _09571_/X _09656_/B1 _18394_/Q vssd1 vssd1 vccd1 vccd1
+ _09572_/X sky130_fd_sc_hd__o32a_1
XFILLER_209_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09006_ _11217_/C _11218_/B _09245_/A vssd1 vssd1 vccd1 vccd1 _09006_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1507 fanout1514/X vssd1 vssd1 vccd1 vccd1 _10224_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1518 fanout1524/X vssd1 vssd1 vccd1 vccd1 _09302_/S sky130_fd_sc_hd__buf_4
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout520 _17219_/Y vssd1 vssd1 vccd1 vccd1 _17244_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_266_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout531 _11729_/X vssd1 vssd1 vccd1 vccd1 _11899_/A sky130_fd_sc_hd__buf_8
Xfanout1529 _10653_/A1 vssd1 vssd1 vccd1 vccd1 _10643_/S sky130_fd_sc_hd__buf_6
Xfanout542 _17540_/B1 vssd1 vssd1 vccd1 vccd1 _15717_/B2 sky130_fd_sc_hd__buf_4
XFILLER_219_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09908_ _09908_/A1 _09907_/A _09907_/B _09908_/B1 _18374_/Q vssd1 vssd1 vccd1 vccd1
+ _09908_/X sky130_fd_sc_hd__o32a_1
XFILLER_263_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout553 _17211_/A vssd1 vssd1 vccd1 vccd1 _17166_/A sky130_fd_sc_hd__buf_4
Xfanout564 _15112_/Y vssd1 vssd1 vccd1 vccd1 _15437_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout575 _16078_/X vssd1 vssd1 vccd1 vccd1 _16096_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_19_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout586 _12088_/A2 vssd1 vssd1 vccd1 vccd1 _12086_/A2 sky130_fd_sc_hd__buf_4
XFILLER_246_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout597 _14268_/B vssd1 vssd1 vccd1 vccd1 _12433_/B sky130_fd_sc_hd__buf_2
X_09839_ _09835_/X _09836_/X _09837_/X _09838_/X _11173_/S _09086_/A vssd1 vssd1 vccd1
+ vccd1 _09839_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12850_ _19234_/Q _13495_/A2 _13495_/B1 _19266_/Q vssd1 vssd1 vccd1 vccd1 _12850_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11801_ _11801_/A _11834_/B vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__nor2_8
XFILLER_262_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _17856_/Q _12919_/A2 _12769_/X _13115_/B2 _12780_/X vssd1 vssd1 vccd1 vccd1
+ _12781_/X sky130_fd_sc_hd__a221o_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _17722_/A0 _18370_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _18370_/D sky130_fd_sc_hd__mux2_1
XFILLER_214_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11732_/A _12900_/A vssd1 vssd1 vccd1 vccd1 _11732_/Y sky130_fd_sc_hd__xnor2_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _18591_/Q _14451_/B vssd1 vssd1 vccd1 vccd1 _18304_/D sky130_fd_sc_hd__and2_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11663_ _11663_/A _11727_/B vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__nor2_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13402_ _13937_/A _13402_/B vssd1 vssd1 vccd1 vccd1 _13402_/X sky130_fd_sc_hd__or2_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10614_ _11584_/A1 _19218_/Q _19186_/Q _10467_/S _11584_/C1 vssd1 vssd1 vccd1 vccd1
+ _10614_/X sky130_fd_sc_hd__a221o_1
X_17170_ _19408_/Q fanout536/X _17473_/A _17120_/B vssd1 vssd1 vccd1 vccd1 _17171_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14382_ _18234_/Q _16490_/A0 _14382_/S vssd1 vssd1 vccd1 vccd1 _18234_/D sky130_fd_sc_hd__mux2_1
XFILLER_195_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11594_ _11594_/A1 _19226_/Q _19194_/Q _11613_/S _08899_/A vssd1 vssd1 vccd1 vccd1
+ _11594_/X sky130_fd_sc_hd__a221o_1
X_16121_ _18763_/Q _16139_/B vssd1 vssd1 vccd1 vccd1 _16121_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13333_ _15380_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _13333_/Y sky130_fd_sc_hd__nand2_1
XFILLER_182_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10545_ _18899_/Q _10838_/B _10544_/X _09095_/A vssd1 vssd1 vccd1 vccd1 _10545_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16052_ _16052_/A _16052_/B vssd1 vssd1 vccd1 vccd1 _18737_/D sky130_fd_sc_hd__and2_1
X_13264_ _13263_/A _12941_/X _13263_/Y _12739_/S vssd1 vssd1 vccd1 vccd1 _13264_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10476_ _10850_/A1 _17783_/Q _10840_/S _18332_/Q vssd1 vssd1 vccd1 vccd1 _10476_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15003_ _15003_/A1 _13954_/Y _15003_/B1 _18657_/Q _15003_/C1 vssd1 vssd1 vccd1 vccd1
+ _15003_/X sky130_fd_sc_hd__a221o_1
X_12215_ _17869_/Q _12216_/C _17870_/Q vssd1 vssd1 vccd1 vccd1 _12217_/B sky130_fd_sc_hd__a21oi_1
X_13195_ _13316_/B _12836_/Y _13195_/S vssd1 vssd1 vccd1 vccd1 _13195_/X sky130_fd_sc_hd__mux2_2
XFILLER_151_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12146_ _17844_/Q _12146_/B vssd1 vssd1 vccd1 vccd1 _12152_/C sky130_fd_sc_hd__and2_2
XFILLER_150_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16954_ _16970_/A1 _17947_/Q _16953_/X vssd1 vssd1 vccd1 vccd1 _17202_/B sky130_fd_sc_hd__o21a_4
XFILLER_111_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12077_ _17816_/Q _12085_/B vssd1 vssd1 vccd1 vccd1 _12077_/X sky130_fd_sc_hd__or2_1
X_15905_ _15905_/A _15905_/B _15905_/C vssd1 vssd1 vccd1 vccd1 _15905_/X sky130_fd_sc_hd__and3_1
XFILLER_265_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11028_ _11511_/A _11028_/B vssd1 vssd1 vccd1 vccd1 _11028_/Y sky130_fd_sc_hd__nand2_1
XFILLER_238_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16885_ _18752_/Q _16893_/A2 _16893_/B1 input216/X _12483_/A vssd1 vssd1 vccd1 vccd1
+ _16885_/X sky130_fd_sc_hd__a221o_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18624_ _19628_/CLK _18624_/D vssd1 vssd1 vccd1 vccd1 _18624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_266_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _18744_/Q _12276_/A _16877_/B1 input237/X vssd1 vssd1 vccd1 vccd1 _15837_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_253_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18555_ _19609_/CLK _18555_/D vssd1 vssd1 vccd1 vccd1 _18555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _15770_/A vssd1 vssd1 vccd1 vccd1 _15767_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12979_ _13929_/A1 _12978_/X _12962_/X vssd1 vssd1 vccd1 vccd1 _12979_/X sky130_fd_sc_hd__a21o_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17506_ _18585_/Q _17544_/A _08883_/A vssd1 vssd1 vccd1 vccd1 _17506_/X sky130_fd_sc_hd__o21a_1
X_14718_ _14718_/A _14718_/B vssd1 vssd1 vccd1 vccd1 _14718_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18486_ _19291_/CLK _18486_/D vssd1 vssd1 vccd1 vccd1 _18486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15698_ _15717_/B2 _15697_/X _15782_/B1 vssd1 vssd1 vccd1 vccd1 _15698_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_480 input231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_491 _18115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17437_ _18110_/Q _17437_/A2 _17435_/X _17436_/X vssd1 vssd1 vccd1 vccd1 _17437_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14649_ _16608_/A0 _18455_/Q _14660_/S vssd1 vssd1 vccd1 vccd1 _18455_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_16 _14909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_27 _17175_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_38 _09139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 _12613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ _17368_/A _17368_/B vssd1 vssd1 vccd1 vccd1 _19481_/D sky130_fd_sc_hd__and2_1
XFILLER_192_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19107_ _19636_/CLK _19107_/D vssd1 vssd1 vccd1 vccd1 _19107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16319_ _17717_/A0 _18932_/Q _16320_/S vssd1 vssd1 vccd1 vccd1 _18932_/D sky130_fd_sc_hd__mux2_1
X_17299_ _18127_/Q _15782_/A1 _17199_/Y _17307_/B vssd1 vssd1 vccd1 vccd1 _17299_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19038_ _19621_/CLK _19038_/D vssd1 vssd1 vccd1 vccd1 _19038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09624_ _10323_/A1 _18138_/Q _18784_/Q _10313_/S _11480_/C1 vssd1 vssd1 vccd1 vccd1
+ _09624_/X sky130_fd_sc_hd__a221o_1
XFILLER_244_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09555_ _10180_/A _09549_/X _09554_/X _09531_/Y _09548_/Y vssd1 vssd1 vccd1 vccd1
+ _09555_/X sky130_fd_sc_hd__a32o_2
Xclkbuf_leaf_37_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19138_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_270_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09486_ input121/X input156/X _09657_/S vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__mux2_8
XFILLER_24_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10330_ _10328_/X _10329_/X _10335_/S vssd1 vssd1 vccd1 vccd1 _10330_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ _09463_/S _10256_/X _10260_/X vssd1 vssd1 vccd1 vccd1 _10261_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_106_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12000_ _17767_/Q _17701_/A0 _12021_/S vssd1 vssd1 vccd1 vccd1 _17767_/D sky130_fd_sc_hd__mux2_1
XFILLER_278_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10192_ _10338_/A1 _10191_/X _11459_/B1 vssd1 vssd1 vccd1 vccd1 _10192_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1304 _12272_/X vssd1 vssd1 vccd1 vccd1 _16893_/A2 sky130_fd_sc_hd__buf_2
Xfanout1315 _12420_/B1 vssd1 vssd1 vccd1 vccd1 _12432_/B1 sky130_fd_sc_hd__buf_6
Xfanout1326 _10260_/B1 vssd1 vssd1 vccd1 vccd1 _11466_/B1 sky130_fd_sc_hd__buf_12
Xfanout1337 _10409_/A vssd1 vssd1 vccd1 vccd1 _09129_/S sky130_fd_sc_hd__buf_6
Xfanout1348 _09919_/C1 vssd1 vssd1 vccd1 vccd1 _09463_/S sky130_fd_sc_hd__buf_6
Xfanout1359 _09093_/Y vssd1 vssd1 vccd1 vccd1 _11224_/B sky130_fd_sc_hd__buf_6
XFILLER_87_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13951_ _19391_/Q _13951_/A2 _13949_/X _13950_/X _13951_/C1 vssd1 vssd1 vccd1 vccd1
+ _13951_/X sky130_fd_sc_hd__o221a_4
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12902_ _11732_/Y _13349_/B _12901_/X _12442_/C vssd1 vssd1 vccd1 vccd1 _12902_/X
+ sky130_fd_sc_hd__a211o_1
X_16670_ _19245_/Q _19244_/Q _16670_/C vssd1 vssd1 vccd1 vccd1 _16673_/B sky130_fd_sc_hd__and3_1
XFILLER_35_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13882_ _19453_/Q _13949_/A2 _13880_/X _13881_/X _13949_/C1 vssd1 vssd1 vccd1 vccd1
+ _13882_/X sky130_fd_sc_hd__o221a_1
XFILLER_207_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15621_ _18585_/Q _18584_/Q _15621_/C vssd1 vssd1 vccd1 vccd1 _15662_/C sky130_fd_sc_hd__and3_2
X_12833_ _12833_/A vssd1 vssd1 vccd1 vccd1 _12833_/Y sky130_fd_sc_hd__inv_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _19618_/CLK _18340_/D vssd1 vssd1 vccd1 vccd1 _18340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15702_/A _15553_/B vssd1 vssd1 vccd1 vccd1 _15580_/A sky130_fd_sc_hd__nor2_2
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12761_/X _13292_/A2 _12763_/X _13256_/B1 _17920_/Q vssd1 vssd1 vccd1 vccd1
+ _12765_/B sky130_fd_sc_hd__a32o_1
XFILLER_226_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14503_ _17705_/A0 _18353_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _18353_/D sky130_fd_sc_hd__mux2_1
X_11715_ _11715_/A _11715_/B _11715_/C _11715_/D vssd1 vssd1 vccd1 vccd1 _14417_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18271_ _18272_/CLK _18271_/D vssd1 vssd1 vccd1 vccd1 _18271_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _15484_/A _15484_/C _15484_/B vssd1 vssd1 vccd1 vccd1 _15486_/A sky130_fd_sc_hd__a21o_1
XFILLER_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12695_ _12694_/X _12693_/X _12818_/S vssd1 vssd1 vccd1 vccd1 _12695_/X sky130_fd_sc_hd__mux2_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17222_ _17220_/Y _17221_/X _14423_/B vssd1 vssd1 vccd1 vccd1 _19424_/D sky130_fd_sc_hd__a21oi_1
X_14434_ _18573_/Q _14451_/B vssd1 vssd1 vccd1 vccd1 _18286_/D sky130_fd_sc_hd__and2_1
X_11646_ _11647_/A _11816_/A vssd1 vssd1 vccd1 vccd1 _11869_/B sky130_fd_sc_hd__nor2_4
XFILLER_156_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 core_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
X_14365_ _18217_/Q _17672_/A0 _14382_/S vssd1 vssd1 vccd1 vccd1 _18217_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput25 core_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_2
X_17153_ _17255_/A _17153_/B vssd1 vssd1 vccd1 vccd1 _19402_/D sky130_fd_sc_hd__nor2_1
X_11577_ _11575_/X _11576_/X _11577_/S vssd1 vssd1 vccd1 vccd1 _11577_/X sky130_fd_sc_hd__mux2_1
Xinput36 core_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_2
Xinput47 dout0[13] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_2
X_16104_ _16142_/A1 _16103_/Y _16149_/A vssd1 vssd1 vccd1 vccd1 _18754_/D sky130_fd_sc_hd__a21oi_1
XFILLER_155_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13316_ _13316_/A _13316_/B vssd1 vssd1 vccd1 vccd1 _13316_/Y sky130_fd_sc_hd__nand2_1
Xinput58 dout0[23] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10528_ _10085_/A _10085_/B _09322_/X _11143_/A1 vssd1 vssd1 vccd1 vccd1 _10528_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17084_ _17589_/A _17108_/A2 _17083_/X _17360_/A vssd1 vssd1 vccd1 vccd1 _19375_/D
+ sky130_fd_sc_hd__o211a_1
Xinput69 dout0[33] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_2
X_14296_ _17714_/A0 _18155_/Q _14301_/S vssd1 vssd1 vccd1 vccd1 _18155_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16035_ _16020_/Y _16034_/X _16033_/X _16052_/A vssd1 vssd1 vccd1 vccd1 _18730_/D
+ sky130_fd_sc_hd__o211a_1
X_13247_ _19370_/Q _13247_/A2 _13245_/X _13246_/X _13247_/C1 vssd1 vssd1 vccd1 vccd1
+ _13247_/X sky130_fd_sc_hd__o221a_4
X_10459_ _17945_/Q _11451_/A2 _10458_/X vssd1 vssd1 vccd1 vccd1 _10459_/X sky130_fd_sc_hd__o21a_4
XFILLER_170_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13178_ _17831_/Q _13105_/B _13176_/X _13177_/X _12548_/X vssd1 vssd1 vccd1 vccd1
+ _13178_/X sky130_fd_sc_hd__o221a_2
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12129_ _12219_/A _12129_/B _12130_/B vssd1 vssd1 vccd1 vccd1 _17837_/D sky130_fd_sc_hd__nor3_1
XFILLER_96_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17986_ _18973_/CLK _17986_/D vssd1 vssd1 vccd1 vccd1 _17986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1860 fanout1863/X vssd1 vssd1 vccd1 vccd1 _14203_/A sky130_fd_sc_hd__clkbuf_2
X_16937_ _18765_/Q _16965_/A2 _16965_/B1 input230/X _16965_/C1 vssd1 vssd1 vccd1 vccd1
+ _16937_/X sky130_fd_sc_hd__a221o_4
Xfanout1871 _17285_/A vssd1 vssd1 vccd1 vccd1 _17210_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1882 _12243_/A vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__buf_4
Xfanout1893 _16737_/A vssd1 vssd1 vccd1 vccd1 _16811_/A sky130_fd_sc_hd__buf_4
XFILLER_265_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16868_ _18748_/Q _12276_/A _16877_/B1 input243/X _08828_/A vssd1 vssd1 vccd1 vccd1
+ _16868_/X sky130_fd_sc_hd__a221o_1
XFILLER_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18607_ _19630_/CLK _18607_/D vssd1 vssd1 vccd1 vccd1 _18607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15819_ _18611_/Q _17709_/A0 _15833_/S vssd1 vssd1 vccd1 vccd1 _18611_/D sky130_fd_sc_hd__mux2_1
X_19587_ _19587_/CLK _19587_/D vssd1 vssd1 vccd1 vccd1 _19587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16799_ _19288_/Q _19287_/Q _16799_/C vssd1 vssd1 vccd1 vccd1 _16802_/B sky130_fd_sc_hd__and3_1
XFILLER_280_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09340_ _10169_/S _09338_/X _09339_/X vssd1 vssd1 vccd1 vccd1 _09340_/X sky130_fd_sc_hd__a21o_1
X_18538_ _18632_/CLK _18538_/D vssd1 vssd1 vccd1 vccd1 _18538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09271_ _09272_/A1 _18213_/Q _09269_/S _18948_/Q _09136_/S vssd1 vssd1 vccd1 vccd1
+ _09271_/X sky130_fd_sc_hd__o221a_1
XFILLER_221_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18469_ _19648_/CLK _18469_/D vssd1 vssd1 vccd1 vccd1 _18469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_155_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19465_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_228_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08986_ _09992_/A _18528_/Q vssd1 vssd1 vccd1 vccd1 _08986_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09607_ _08904_/A _09601_/X _09604_/X _09606_/X _11495_/B1 vssd1 vssd1 vccd1 vccd1
+ _09608_/B sky130_fd_sc_hd__a311o_1
XFILLER_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09538_ _12468_/B _18139_/Q _18785_/Q _09925_/S _09457_/A vssd1 vssd1 vccd1 vccd1
+ _09538_/X sky130_fd_sc_hd__a221o_1
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09469_ _09448_/X _09451_/X _09468_/X vssd1 vssd1 vccd1 vccd1 _09469_/X sky130_fd_sc_hd__a21o_1
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11500_ _18855_/Q _18887_/Q _19047_/Q _19015_/Q _09966_/S _11503_/S1 vssd1 vssd1
+ vccd1 vccd1 _11500_/X sky130_fd_sc_hd__mux4_1
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12480_ _16852_/A _08841_/Y _12478_/Y vssd1 vssd1 vccd1 vccd1 _12554_/A sky130_fd_sc_hd__a21o_1
XFILLER_185_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ _11431_/A _11431_/B vssd1 vssd1 vccd1 vccd1 _11431_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14150_ _14150_/A _14150_/B vssd1 vssd1 vccd1 vccd1 _14151_/D sky130_fd_sc_hd__or2_2
XFILLER_256_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11362_ _11606_/S _11361_/X _11608_/C1 vssd1 vssd1 vccd1 vccd1 _11362_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13101_ _15238_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13101_/Y sky130_fd_sc_hd__nand2_1
X_10313_ _19645_/Q _18934_/Q _10313_/S vssd1 vssd1 vccd1 vccd1 _10313_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14081_ _16597_/A0 _18021_/Q _14104_/S vssd1 vssd1 vccd1 vccd1 _18021_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11293_ _11293_/A _11293_/B vssd1 vssd1 vccd1 vccd1 _12626_/A sky130_fd_sc_hd__nor2_4
XFILLER_152_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _13033_/A _13033_/B vssd1 vssd1 vccd1 vccd1 _13032_/Y sky130_fd_sc_hd__nor2_1
X_10244_ _10263_/A1 _19223_/Q _19191_/Q _10253_/C _11397_/A1 vssd1 vssd1 vccd1 vccd1
+ _10244_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1101 _08882_/Y vssd1 vssd1 vccd1 vccd1 _17426_/B1 sky130_fd_sc_hd__buf_2
XFILLER_279_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17840_ _19310_/CLK _17840_/D vssd1 vssd1 vccd1 vccd1 _17840_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1112 _13637_/A vssd1 vssd1 vccd1 vccd1 _13757_/A sky130_fd_sc_hd__buf_4
X_10175_ _10173_/X _10174_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _10175_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1123 _13791_/A vssd1 vssd1 vccd1 vccd1 _13079_/A sky130_fd_sc_hd__buf_2
XFILLER_239_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1134 _13970_/B2 vssd1 vssd1 vccd1 vccd1 _13936_/B2 sky130_fd_sc_hd__buf_4
XFILLER_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1145 _10194_/C1 vssd1 vssd1 vccd1 vccd1 _10239_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1156 _16004_/C1 vssd1 vssd1 vccd1 vccd1 _16018_/C1 sky130_fd_sc_hd__buf_4
X_17771_ _19599_/CLK _17771_/D vssd1 vssd1 vccd1 vccd1 _17771_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1167 _15851_/Y vssd1 vssd1 vccd1 vccd1 _15906_/B1 sky130_fd_sc_hd__buf_4
X_14983_ _14992_/A1 _13886_/X _14983_/B1 _18655_/Q _14741_/B vssd1 vssd1 vccd1 vccd1
+ _14983_/X sky130_fd_sc_hd__a221o_1
XFILLER_281_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1178 _13260_/Y vssd1 vssd1 vccd1 vccd1 _13909_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1189 _08946_/Y vssd1 vssd1 vccd1 vccd1 _08948_/B sky130_fd_sc_hd__buf_8
X_19510_ _19519_/CLK _19510_/D vssd1 vssd1 vccd1 vccd1 _19510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16722_ _19260_/Q _19259_/Q _16722_/C vssd1 vssd1 vccd1 vccd1 _16728_/C sky130_fd_sc_hd__and3_1
X_13934_ _18131_/Q _13934_/B vssd1 vssd1 vccd1 vccd1 _13935_/B sky130_fd_sc_hd__or2_1
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19441_ _19507_/CLK _19441_/D vssd1 vssd1 vccd1 vccd1 _19441_/Q sky130_fd_sc_hd__dfxtp_1
X_16653_ _19238_/Q _19237_/Q _19234_/Q _16653_/D vssd1 vssd1 vccd1 vccd1 _16677_/B
+ sky130_fd_sc_hd__and4_1
X_13865_ _13259_/X _13859_/X _13861_/Y _13864_/X vssd1 vssd1 vccd1 vccd1 _13865_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_263_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15604_ _18584_/Q _15621_/C vssd1 vssd1 vccd1 vccd1 _15604_/X sky130_fd_sc_hd__or2_1
XFILLER_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19372_ _19502_/CLK _19372_/D vssd1 vssd1 vccd1 vccd1 _19372_/Q sky130_fd_sc_hd__dfxtp_1
X_12816_ _12811_/X _12815_/Y _13041_/S vssd1 vssd1 vccd1 vccd1 _12817_/A sky130_fd_sc_hd__mux2_1
X_16584_ _16617_/A0 _19188_/Q _16585_/S vssd1 vssd1 vccd1 vccd1 _19188_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13796_ _13807_/B _13961_/A _13795_/X vssd1 vssd1 vccd1 vccd1 _13796_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18323_ _19602_/CLK _18323_/D vssd1 vssd1 vccd1 vccd1 _18323_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ _15581_/C _15535_/B vssd1 vssd1 vccd1 vccd1 _15538_/B sky130_fd_sc_hd__nor2_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12747_ _12813_/S _13958_/B _12707_/X vssd1 vssd1 vccd1 vccd1 _12748_/A sky130_fd_sc_hd__o21ai_2
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _19075_/CLK _18254_/D vssd1 vssd1 vccd1 vccd1 _18254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12678_ _12677_/X _12676_/X _12823_/A vssd1 vssd1 vccd1 vccd1 _12678_/X sky130_fd_sc_hd__mux2_1
X_15466_ _18577_/Q _15465_/C _18578_/Q vssd1 vssd1 vccd1 vccd1 _15467_/B sky130_fd_sc_hd__a21oi_1
XFILLER_175_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17205_ _17208_/A _17205_/B vssd1 vssd1 vccd1 vccd1 _17205_/Y sky130_fd_sc_hd__nand2_1
X_14417_ _14417_/A _14417_/B _14417_/C vssd1 vssd1 vccd1 vccd1 _18274_/D sky130_fd_sc_hd__and3_4
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11629_ _11627_/Y _11629_/B vssd1 vssd1 vccd1 vccd1 _12656_/B sky130_fd_sc_hd__and2b_4
X_18185_ _19219_/CLK _18185_/D vssd1 vssd1 vccd1 vccd1 _18185_/Q sky130_fd_sc_hd__dfxtp_1
X_15397_ _19469_/Q _19403_/Q vssd1 vssd1 vccd1 vccd1 _15398_/B sky130_fd_sc_hd__or2_1
XFILLER_129_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17136_ _17157_/A _17569_/A vssd1 vssd1 vccd1 vccd1 _17418_/A sky130_fd_sc_hd__nand2_1
XFILLER_184_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14348_ _17533_/A _17210_/A vssd1 vssd1 vccd1 vccd1 _18303_/D sky130_fd_sc_hd__nor2_1
XFILLER_128_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14279_ _16597_/A0 _18138_/Q _14301_/S vssd1 vssd1 vccd1 vccd1 _18138_/D sky130_fd_sc_hd__mux2_1
X_17067_ _19367_/Q _17077_/B vssd1 vssd1 vccd1 vccd1 _17067_/X sky130_fd_sc_hd__or2_1
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16018_ _18724_/Q _15953_/B _16147_/A2 _18773_/Q _16018_/C1 vssd1 vssd1 vccd1 vccd1
+ _16018_/X sky130_fd_sc_hd__a221o_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _17915_/Q vssd1 vssd1 vccd1 vccd1 _08840_/Y sky130_fd_sc_hd__inv_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17969_ _17975_/CLK _17969_/D vssd1 vssd1 vccd1 vccd1 _17969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1690 _08845_/Y vssd1 vssd1 vccd1 vccd1 _12468_/B sky130_fd_sc_hd__buf_8
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19639_ _19639_/CLK _19639_/D vssd1 vssd1 vccd1 vccd1 _19639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09323_ input114/X input149/X _09657_/S vssd1 vssd1 vccd1 vccd1 _09323_/X sky130_fd_sc_hd__mux2_8
XFILLER_179_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09254_ _10409_/A _09252_/X _09253_/X vssd1 vssd1 vccd1 vccd1 _09254_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09185_ _10336_/A _09183_/X _09184_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09186_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_175_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput204 localMemory_wb_adr_i[22] vssd1 vssd1 vccd1 vccd1 _12269_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_216_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput215 localMemory_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input215/X sky130_fd_sc_hd__clkbuf_16
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput226 localMemory_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input226/X sky130_fd_sc_hd__clkbuf_16
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 localMemory_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input237/X sky130_fd_sc_hd__clkbuf_16
XFILLER_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19628_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput248 localMemory_wb_sel_i[1] vssd1 vssd1 vccd1 vccd1 input248/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput259 manufacturerID[5] vssd1 vssd1 vccd1 vccd1 _15872_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_276_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08969_ _09976_/A1 _08968_/X _11515_/B1 vssd1 vssd1 vccd1 vccd1 _08969_/X sky130_fd_sc_hd__a21o_1
XFILLER_236_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ _18693_/Q _11977_/B _11977_/X vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__a21bo_1
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10931_ _19054_/Q _19022_/Q _10940_/S vssd1 vssd1 vccd1 vccd1 _10931_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13650_ _19254_/Q _13943_/A2 _13943_/B1 _19286_/Q vssd1 vssd1 vccd1 vccd1 _13650_/X
+ sky130_fd_sc_hd__a22o_2
X_10862_ _11312_/A1 _18614_/Q _18185_/Q _10864_/S vssd1 vssd1 vccd1 vccd1 _10862_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12601_ _13263_/A _12601_/B vssd1 vssd1 vccd1 vccd1 _12601_/Y sky130_fd_sc_hd__nand2_1
XFILLER_231_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _13581_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13581_/X sky130_fd_sc_hd__or2_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10793_ _11103_/A _11860_/A vssd1 vssd1 vccd1 vccd1 _10793_/Y sky130_fd_sc_hd__nor2_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ _13165_/B _13165_/C vssd1 vssd1 vccd1 vccd1 _12532_/Y sky130_fd_sc_hd__nor2_2
XFILLER_169_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15320_ _19466_/Q _19400_/Q vssd1 vssd1 vccd1 vccd1 _15321_/B sky130_fd_sc_hd__nand2_1
XFILLER_223_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12463_ _16852_/A _14004_/A _14992_/A1 vssd1 vssd1 vccd1 vccd1 _12463_/X sky130_fd_sc_hd__a21o_4
X_15251_ _19431_/Q _15411_/B _17151_/A _15250_/X vssd1 vssd1 vccd1 vccd1 _15251_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11414_ _11512_/A1 _19599_/Q _19567_/Q _11426_/B2 vssd1 vssd1 vccd1 vccd1 _11414_/X
+ sky130_fd_sc_hd__a22o_1
X_14202_ _18712_/Q _18099_/Q _14204_/S vssd1 vssd1 vccd1 vccd1 _14203_/B sky130_fd_sc_hd__mux2_1
XFILLER_172_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15182_ _18565_/Q _18564_/Q _18566_/Q vssd1 vssd1 vccd1 vccd1 _15183_/B sky130_fd_sc_hd__a21oi_1
X_12394_ _12408_/B _12394_/B vssd1 vssd1 vccd1 vccd1 _12394_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14133_ _10532_/B _18072_/Q _14140_/S vssd1 vssd1 vccd1 vccd1 _18072_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11345_ _11360_/A1 _18147_/Q _18793_/Q _11360_/B2 vssd1 vssd1 vccd1 vccd1 _11345_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14064_ _17681_/A0 _18006_/Q _14064_/S vssd1 vssd1 vccd1 vccd1 _18006_/D sky130_fd_sc_hd__mux2_1
X_18941_ _19133_/CLK _18941_/D vssd1 vssd1 vccd1 vccd1 _18941_/Q sky130_fd_sc_hd__dfxtp_1
X_11276_ _11277_/A1 _18954_/Q _18219_/Q _11284_/B2 vssd1 vssd1 vccd1 vccd1 _11276_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13015_ _19495_/Q _13064_/B _13243_/B1 _13014_/X vssd1 vssd1 vccd1 vccd1 _13015_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_279_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10227_ _08896_/A _10226_/X _11501_/B1 vssd1 vssd1 vccd1 vccd1 _10227_/X sky130_fd_sc_hd__a21o_1
X_18872_ _19193_/CLK _18872_/D vssd1 vssd1 vccd1 vccd1 _18872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_279_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17823_ _18761_/CLK _17823_/D vssd1 vssd1 vccd1 vccd1 _17823_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10158_ _10159_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__and2_2
XFILLER_282_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17754_ _18654_/Q vssd1 vssd1 vccd1 vccd1 _18654_/D sky130_fd_sc_hd__clkbuf_2
X_10089_ _11452_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10089_/Y sky130_fd_sc_hd__nor2_1
X_14966_ _14996_/A1 _14965_/X _15006_/B1 vssd1 vssd1 vccd1 vccd1 _14966_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_48_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16705_ _16795_/A _16705_/B _16706_/B vssd1 vssd1 vccd1 vccd1 _19254_/D sky130_fd_sc_hd__nor3_1
XFILLER_75_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13917_ _13917_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _13917_/Y sky130_fd_sc_hd__nor2_1
X_17685_ _17685_/A0 _19612_/Q _17689_/S vssd1 vssd1 vccd1 vccd1 _19612_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14897_ _14897_/A vssd1 vssd1 vccd1 vccd1 _14897_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19424_ _19526_/CLK _19424_/D vssd1 vssd1 vccd1 vccd1 _19424_/Q sky130_fd_sc_hd__dfxtp_1
X_16636_ _19234_/Q _16677_/A _16635_/Y vssd1 vssd1 vccd1 vccd1 _19234_/D sky130_fd_sc_hd__o21a_1
XFILLER_251_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13848_ _19550_/Q _13946_/B vssd1 vssd1 vccd1 vccd1 _13848_/X sky130_fd_sc_hd__or2_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19355_ _19483_/CLK _19355_/D vssd1 vssd1 vccd1 vccd1 _19355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16567_ _17700_/A0 _19171_/Q _16589_/S vssd1 vssd1 vccd1 vccd1 _19171_/D sky130_fd_sc_hd__mux2_1
X_13779_ _17881_/Q _13847_/A2 _13777_/X _13928_/A1 _13854_/B1 vssd1 vssd1 vccd1 vccd1
+ _13779_/X sky130_fd_sc_hd__a221o_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18306_ _19444_/CLK _18306_/D vssd1 vssd1 vccd1 vccd1 _18306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15518_ _15497_/A _15496_/B _15496_/A vssd1 vssd1 vccd1 vccd1 _15522_/A sky130_fd_sc_hd__a21boi_4
X_19286_ _19286_/CLK _19286_/D vssd1 vssd1 vccd1 vccd1 _19286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16498_ _17664_/A0 _19104_/Q _16515_/S vssd1 vssd1 vccd1 vccd1 _19104_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ _19619_/CLK _18237_/D vssd1 vssd1 vccd1 vccd1 _18237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15449_ _10513_/S _15452_/A _15484_/A vssd1 vssd1 vccd1 vccd1 _15455_/A sky130_fd_sc_hd__o21a_1
XFILLER_191_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18168_ _19148_/CLK _18168_/D vssd1 vssd1 vccd1 vccd1 _18168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17119_ _17199_/A _17119_/B vssd1 vssd1 vccd1 vccd1 _17119_/X sky130_fd_sc_hd__and2_1
X_18099_ _18715_/CLK _18099_/D vssd1 vssd1 vccd1 vccd1 _18099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09941_ _10180_/A _09940_/X _09924_/X _11024_/A1 vssd1 vssd1 vccd1 vccd1 _09941_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout905 _16454_/S vssd1 vssd1 vccd1 vccd1 _16457_/S sky130_fd_sc_hd__buf_12
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout916 _16278_/S vssd1 vssd1 vccd1 vccd1 _16292_/S sky130_fd_sc_hd__buf_12
Xfanout927 _16194_/X vssd1 vssd1 vccd1 vccd1 _16212_/S sky130_fd_sc_hd__buf_12
XFILLER_258_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _18238_/Q _18813_/Q _18441_/Q _18342_/Q _10054_/S _08874_/D vssd1 vssd1 vccd1
+ vccd1 _09872_/X sky130_fd_sc_hd__mux4_1
Xfanout938 _14673_/X vssd1 vssd1 vccd1 vccd1 _14982_/B sky130_fd_sc_hd__buf_4
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout949 _14648_/S vssd1 vssd1 vccd1 vccd1 _14664_/S sky130_fd_sc_hd__buf_12
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08823_ _18777_/Q vssd1 vssd1 vccd1 vccd1 _14423_/A sky130_fd_sc_hd__inv_2
XFILLER_273_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_7__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_258_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_309 _18113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_170_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19450_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09306_ _19076_/Q _18980_/Q _09306_/S vssd1 vssd1 vccd1 vccd1 _09306_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09237_ _18390_/Q _09656_/B1 _09236_/Y _09992_/A vssd1 vssd1 vccd1 vccd1 _09901_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_166_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09168_ _19045_/Q _19013_/Q _10099_/S vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09099_ _09099_/A _09285_/C vssd1 vssd1 vccd1 vccd1 _09099_/Y sky130_fd_sc_hd__nand2_8
X_11130_ _11106_/Y _11110_/Y _11621_/C1 vssd1 vssd1 vccd1 vccd1 _11130_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11061_ _12594_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11062_/B sky130_fd_sc_hd__nor2_4
XFILLER_122_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10012_ _10010_/X _10011_/X _10707_/A vssd1 vssd1 vccd1 vccd1 _10012_/X sky130_fd_sc_hd__mux2_1
XFILLER_276_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _12051_/A _14819_/X _14993_/S vssd1 vssd1 vccd1 vccd1 _14820_/X sky130_fd_sc_hd__mux2_1
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _14912_/A1 _13076_/Y _14973_/B1 _18632_/Q _14741_/B vssd1 vssd1 vccd1 vccd1
+ _14751_/X sky130_fd_sc_hd__a221o_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11963_ _18509_/Q _11720_/X _11913_/X _11706_/X vssd1 vssd1 vccd1 vccd1 _11963_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _13259_/X _13695_/X _13698_/Y _13701_/X vssd1 vssd1 vccd1 vccd1 _13702_/X
+ sky130_fd_sc_hd__a31o_1
X_17470_ _13476_/B _17520_/A2 _17532_/A2 _17806_/Q _17550_/A vssd1 vssd1 vccd1 vccd1
+ _17470_/X sky130_fd_sc_hd__a221o_1
X_10914_ _18990_/Q _11300_/B vssd1 vssd1 vccd1 vccd1 _10914_/X sky130_fd_sc_hd__or2_1
XFILLER_232_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _14682_/A _14688_/C vssd1 vssd1 vccd1 vccd1 _14683_/B sky130_fd_sc_hd__nor2_2
X_11894_ _11899_/A _11894_/B _11894_/C vssd1 vssd1 vccd1 vccd1 _11894_/X sky130_fd_sc_hd__and3_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16421_ _16619_/A0 _19030_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _19030_/D sky130_fd_sc_hd__mux2_1
XFILLER_260_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10845_ _18552_/Q _10853_/S vssd1 vssd1 vccd1 vccd1 _10845_/X sky130_fd_sc_hd__or2_1
XFILLER_60_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13633_ _19381_/Q _13951_/A2 _13631_/X _13632_/X _13951_/C1 vssd1 vssd1 vccd1 vccd1
+ _13633_/X sky130_fd_sc_hd__o221a_4
XFILLER_232_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19140_ _19140_/CLK _19140_/D vssd1 vssd1 vccd1 vccd1 _19140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16352_ _18964_/Q _16551_/A0 _16352_/S vssd1 vssd1 vccd1 vccd1 _18964_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10776_ _18553_/Q _18428_/Q _18037_/Q _18005_/Q _10853_/S _11311_/C1 vssd1 vssd1
+ vccd1 vccd1 _10776_/X sky130_fd_sc_hd__mux4_1
X_13564_ _13462_/A _13562_/Y _13563_/X _12448_/D _15426_/B vssd1 vssd1 vccd1 vccd1
+ _13564_/X sky130_fd_sc_hd__a311o_2
XFILLER_157_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15303_ _15303_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _15303_/X sky130_fd_sc_hd__and2_1
XFILLER_200_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12515_ _12577_/A _12552_/A vssd1 vssd1 vccd1 vccd1 _12584_/A sky130_fd_sc_hd__or2_4
X_19071_ _19634_/CLK _19071_/D vssd1 vssd1 vccd1 vccd1 _19071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13495_ _19249_/Q _13495_/A2 _13495_/B1 _19281_/Q vssd1 vssd1 vccd1 vccd1 _13495_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_201_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16283_ _17714_/A0 _18897_/Q _16288_/S vssd1 vssd1 vccd1 vccd1 _18897_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18022_ _18445_/CLK _18022_/D vssd1 vssd1 vccd1 vccd1 _18022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12446_ _12442_/B _12443_/B _09068_/C _12438_/B vssd1 vssd1 vccd1 vccd1 _12446_/X
+ sky130_fd_sc_hd__a211o_1
X_15234_ _19462_/Q _15233_/Y _15400_/S vssd1 vssd1 vccd1 vccd1 _15234_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ _17900_/Q _12408_/B _12376_/Y _13981_/C1 vssd1 vssd1 vccd1 vccd1 _17900_/D
+ sky130_fd_sc_hd__o211a_1
X_15165_ _19459_/Q _19393_/Q vssd1 vssd1 vccd1 vccd1 _15166_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14116_ _16500_/A0 _18055_/Q _14137_/S vssd1 vssd1 vccd1 vccd1 _18055_/D sky130_fd_sc_hd__mux2_1
X_11328_ _11324_/X _11327_/X _11328_/S vssd1 vssd1 vccd1 vccd1 _11328_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15096_ _19384_/Q _15086_/B input185/X _15088_/X vssd1 vssd1 vccd1 vccd1 _15096_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18924_ _19635_/CLK _18924_/D vssd1 vssd1 vccd1 vccd1 _18924_/Q sky130_fd_sc_hd__dfxtp_1
X_14047_ _16597_/A0 _17989_/Q _14070_/S vssd1 vssd1 vccd1 vccd1 _17989_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11259_ _09494_/A _11490_/B _11489_/B1 _11258_/Y vssd1 vssd1 vccd1 vccd1 _12595_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_262_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18855_ _19627_/CLK _18855_/D vssd1 vssd1 vccd1 vccd1 _18855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17806_ _17814_/CLK _17806_/D vssd1 vssd1 vccd1 vccd1 _17806_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18786_ _18880_/CLK _18786_/D vssd1 vssd1 vccd1 vccd1 _18786_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ _18714_/Q _16002_/A2 _16004_/B1 _18763_/Q _16004_/C1 vssd1 vssd1 vccd1 vccd1
+ _15998_/X sky130_fd_sc_hd__a221o_1
XFILLER_209_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17737_ _18637_/Q vssd1 vssd1 vccd1 vccd1 _18637_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_282_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ _14979_/A1 _18272_/Q _14948_/Y _11712_/A vssd1 vssd1 vccd1 vccd1 _14949_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17668_ _17668_/A0 _19595_/Q _17687_/S vssd1 vssd1 vccd1 vccd1 _19595_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19407_ _19543_/CLK _19407_/D vssd1 vssd1 vccd1 vccd1 _19407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16619_ _16619_/A0 _19222_/Q _16619_/S vssd1 vssd1 vccd1 vccd1 _19222_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17599_ _19488_/Q _15092_/X _17556_/A _17178_/B _17556_/X vssd1 vssd1 vccd1 vccd1
+ _17599_/X sky130_fd_sc_hd__a221o_1
XFILLER_250_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19338_ _19399_/CLK _19338_/D vssd1 vssd1 vccd1 vccd1 _19338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19269_ _19273_/CLK _19269_/D vssd1 vssd1 vccd1 vccd1 _19269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09022_ _09043_/A _09009_/X _09028_/B vssd1 vssd1 vccd1 vccd1 _09022_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout702 _12544_/Y vssd1 vssd1 vccd1 vccd1 _13625_/A2 sky130_fd_sc_hd__buf_2
X_09924_ _09922_/X _09923_/X _09089_/Y vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__o21a_1
Xfanout713 _12919_/A2 vssd1 vssd1 vccd1 vccd1 _13747_/A2 sky130_fd_sc_hd__buf_4
XFILLER_277_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout724 _12495_/Y vssd1 vssd1 vccd1 vccd1 _13744_/A2 sky130_fd_sc_hd__buf_4
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout735 _11375_/X vssd1 vssd1 vccd1 vccd1 _11376_/B sky130_fd_sc_hd__buf_4
Xfanout746 _13314_/S vssd1 vssd1 vccd1 vccd1 _13135_/S sky130_fd_sc_hd__buf_4
XFILLER_274_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout757 _17702_/A0 vssd1 vssd1 vccd1 vccd1 _16602_/A0 sky130_fd_sc_hd__clkbuf_4
X_09855_ _19588_/Q _10001_/S _09853_/S _09854_/X vssd1 vssd1 vccd1 vccd1 _09855_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_259_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout768 _17691_/Y vssd1 vssd1 vccd1 vccd1 _17723_/S sky130_fd_sc_hd__buf_12
XFILLER_58_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout779 _16623_/S vssd1 vssd1 vccd1 vccd1 _16619_/S sky130_fd_sc_hd__buf_12
XFILLER_283_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09786_ _18846_/Q _18878_/Q _09797_/S vssd1 vssd1 vccd1 vccd1 _09786_/X sky130_fd_sc_hd__mux2_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_106 _11719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_128 _11806_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _11836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10630_ _10850_/A1 _18227_/Q _10634_/S0 _18962_/Q vssd1 vssd1 vccd1 vccd1 _10630_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_197_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10561_ _10558_/X _10560_/X _10399_/A vssd1 vssd1 vccd1 vccd1 _10561_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_195_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12300_ _18504_/Q _18505_/Q _12277_/B _12299_/X vssd1 vssd1 vccd1 vccd1 _12301_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13280_ _19467_/Q _12529_/Y _12578_/Y _19339_/Q _13279_/X vssd1 vssd1 vccd1 vccd1
+ _13280_/X sky130_fd_sc_hd__a221o_1
XFILLER_212_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10492_ _18557_/Q _18432_/Q _10500_/S vssd1 vssd1 vccd1 vccd1 _10492_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ _17875_/Q _12232_/C _17876_/Q vssd1 vssd1 vccd1 vccd1 _12233_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12162_ _17850_/Q _12162_/B vssd1 vssd1 vccd1 vccd1 _12168_/C sky130_fd_sc_hd__and2_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11113_ _11284_/A1 _18956_/Q _18221_/Q _11125_/B2 vssd1 vssd1 vccd1 vccd1 _11113_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12093_ _17823_/Q _17824_/Q _12092_/Y vssd1 vssd1 vccd1 vccd1 _17824_/D sky130_fd_sc_hd__o21a_1
X_16970_ _16970_/A1 _17951_/Q _16969_/X vssd1 vssd1 vccd1 vccd1 _17214_/B sky130_fd_sc_hd__o21a_4
XFILLER_111_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15921_ _18682_/Q _15948_/A2 _15948_/C1 _15920_/X vssd1 vssd1 vccd1 vccd1 _15921_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ _09967_/S _11043_/X _11501_/B1 vssd1 vssd1 vccd1 vccd1 _11044_/X sky130_fd_sc_hd__a21o_1
XFILLER_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ _19586_/CLK _18640_/D vssd1 vssd1 vccd1 vccd1 _18640_/Q sky130_fd_sc_hd__dfxtp_4
X_15852_ _15853_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15852_/X sky130_fd_sc_hd__and2_2
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _14875_/A1 _14802_/X _14875_/B1 vssd1 vssd1 vccd1 vccd1 _14803_/Y sky130_fd_sc_hd__o21ai_2
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _19433_/CLK _18571_/D vssd1 vssd1 vccd1 vccd1 _18571_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _18592_/Q _15800_/A2 _15775_/X _15782_/X _17376_/A vssd1 vssd1 vccd1 vccd1
+ _18592_/D sky130_fd_sc_hd__o221a_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12995_ _12675_/X _12699_/X _13130_/A vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__mux2_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17522_ _18127_/Q _17539_/C1 _17214_/A _17199_/B vssd1 vssd1 vccd1 vccd1 _17522_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _14732_/X _14733_/X _14995_/A1 vssd1 vssd1 vccd1 vccd1 _14734_/X sky130_fd_sc_hd__a21o_1
XFILLER_18_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _11953_/B2 _11886_/B _11886_/C _11953_/A2 input233/X vssd1 vssd1 vccd1 vccd1
+ _11946_/X sky130_fd_sc_hd__a32o_4
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17453_ _17453_/A _17453_/B vssd1 vssd1 vccd1 vccd1 _17453_/Y sky130_fd_sc_hd__nand2_1
X_14665_ _15835_/B _12277_/B _11719_/X vssd1 vssd1 vccd1 vccd1 _14665_/X sky130_fd_sc_hd__a21bo_1
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11877_ _11803_/Y _11875_/Y _11876_/X vssd1 vssd1 vccd1 vccd1 _11878_/C sky130_fd_sc_hd__o21ai_2
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16404_ _16602_/A0 _19013_/Q _16424_/S vssd1 vssd1 vccd1 vccd1 _19013_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13616_ _13616_/A _13616_/B vssd1 vssd1 vccd1 vccd1 _14149_/A sky130_fd_sc_hd__xnor2_1
XFILLER_60_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10828_ _13623_/A vssd1 vssd1 vccd1 vccd1 _10828_/Y sky130_fd_sc_hd__inv_2
X_17384_ _19488_/Q _17386_/B _17383_/X vssd1 vssd1 vccd1 vccd1 _17384_/X sky130_fd_sc_hd__a21o_1
X_14596_ _14596_/A _14596_/B vssd1 vssd1 vccd1 vccd1 _18405_/D sky130_fd_sc_hd__nor2_1
X_19123_ _19155_/CLK _19123_/D vssd1 vssd1 vccd1 vccd1 _19123_/Q sky130_fd_sc_hd__dfxtp_1
X_16335_ _18947_/Q _16501_/A0 _16357_/S vssd1 vssd1 vccd1 vccd1 _18947_/D sky130_fd_sc_hd__mux2_1
X_13547_ _17938_/Q _13940_/A2 _13546_/X _14181_/A vssd1 vssd1 vccd1 vccd1 _17938_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10759_ _11143_/A1 _10757_/Y _10758_/X vssd1 vssd1 vccd1 vccd1 _10759_/X sky130_fd_sc_hd__o21a_1
XFILLER_146_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19054_ _19632_/CLK _19054_/D vssd1 vssd1 vccd1 vccd1 _19054_/Q sky130_fd_sc_hd__dfxtp_1
X_16266_ _16597_/A0 _18880_/Q _16288_/S vssd1 vssd1 vccd1 vccd1 _18880_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13478_ _17936_/Q _13742_/A2 _13477_/X _14177_/A vssd1 vssd1 vccd1 vccd1 _17936_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18005_ _19600_/CLK _18005_/D vssd1 vssd1 vccd1 vccd1 _18005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15217_ _12318_/A _15215_/Y _15216_/X vssd1 vssd1 vccd1 vccd1 _15219_/B sky130_fd_sc_hd__o21a_2
X_12429_ _12429_/A1 _09232_/A _09484_/X _12429_/B1 _18403_/Q vssd1 vssd1 vccd1 vccd1
+ _12430_/B sky130_fd_sc_hd__o32ai_4
XFILLER_142_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput305 _11725_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[0] sky130_fd_sc_hd__buf_4
X_16197_ _17661_/A0 _18813_/Q _16212_/S vssd1 vssd1 vccd1 vccd1 _18813_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput316 _11726_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[1] sky130_fd_sc_hd__buf_4
Xoutput327 _11738_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[4] sky130_fd_sc_hd__buf_4
Xoutput338 _11827_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[13] sky130_fd_sc_hd__buf_4
X_15148_ _18564_/Q _15351_/A2 _15147_/Y vssd1 vssd1 vccd1 vccd1 _18564_/D sky130_fd_sc_hd__o21a_1
Xoutput349 _11872_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[23] sky130_fd_sc_hd__buf_4
XFILLER_259_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15079_ _18563_/Q _17690_/A0 _15079_/S vssd1 vssd1 vccd1 vccd1 _18563_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18907_ _19618_/CLK _18907_/D vssd1 vssd1 vccd1 vccd1 _18907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_268_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09640_ _09690_/A _09633_/Y _09639_/Y _09350_/S vssd1 vssd1 vccd1 vccd1 _09640_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18838_ _18902_/CLK _18838_/D vssd1 vssd1 vccd1 vccd1 _18838_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_109_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19268_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09571_ input120/X input155/X _09657_/S vssd1 vssd1 vccd1 vccd1 _09571_/X sky130_fd_sc_hd__mux2_8
XFILLER_243_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18769_ _18772_/CLK _18769_/D vssd1 vssd1 vccd1 vccd1 _18769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_283_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09005_ _11691_/B1 _12432_/A2 _09004_/X _09650_/B1 _18404_/Q vssd1 vssd1 vccd1 vccd1
+ _11218_/B sky130_fd_sc_hd__o32a_2
XFILLER_247_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout510 _17423_/B vssd1 vssd1 vccd1 vccd1 _17453_/B sky130_fd_sc_hd__buf_4
XFILLER_59_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1508 fanout1514/X vssd1 vssd1 vccd1 vccd1 _10141_/S sky130_fd_sc_hd__buf_6
Xfanout1519 _11513_/B2 vssd1 vssd1 vccd1 vccd1 _11426_/B2 sky130_fd_sc_hd__buf_6
Xfanout521 _15718_/A2 vssd1 vssd1 vccd1 vccd1 _15800_/A2 sky130_fd_sc_hd__buf_6
XFILLER_120_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09907_ _09907_/A _09907_/B vssd1 vssd1 vccd1 vccd1 _09907_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout532 _11664_/X vssd1 vssd1 vccd1 vccd1 _11706_/B sky130_fd_sc_hd__buf_8
XFILLER_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout543 _15476_/A1 vssd1 vssd1 vccd1 vccd1 _17540_/B1 sky130_fd_sc_hd__buf_6
Xfanout554 _15122_/Y vssd1 vssd1 vccd1 vccd1 _17211_/A sky130_fd_sc_hd__buf_6
XFILLER_259_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout565 _15786_/A2 vssd1 vssd1 vccd1 vccd1 _15763_/A2 sky130_fd_sc_hd__buf_4
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout576 _12379_/A vssd1 vssd1 vccd1 vccd1 _12382_/A sky130_fd_sc_hd__buf_4
XFILLER_86_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout587 _12024_/Y vssd1 vssd1 vccd1 vccd1 _12088_/A2 sky130_fd_sc_hd__buf_4
X_09838_ _11157_/A1 _18135_/Q _18781_/Q _11147_/S vssd1 vssd1 vccd1 vccd1 _09838_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout598 _11697_/Y vssd1 vssd1 vccd1 vccd1 _14268_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09769_ _18442_/Q _18343_/Q _09770_/S vssd1 vssd1 vccd1 vccd1 _09769_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _15082_/B _11800_/B _11800_/C _11800_/D vssd1 vssd1 vccd1 vccd1 _11834_/B
+ sky130_fd_sc_hd__nand4_4
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12779_/X _15860_/A _12918_/S vssd1 vssd1 vccd1 vccd1 _12780_/X sky130_fd_sc_hd__mux2_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11731_ _09897_/Y _11731_/B vssd1 vssd1 vccd1 vccd1 _12900_/A sky130_fd_sc_hd__and2b_4
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _18589_/Q _14450_/B vssd1 vssd1 vccd1 vccd1 _18302_/D sky130_fd_sc_hd__and2_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _15082_/B _15120_/B vssd1 vssd1 vccd1 vccd1 _11727_/B sky130_fd_sc_hd__nand2_4
XFILLER_109_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ _13937_/A _13401_/B vssd1 vssd1 vccd1 vccd1 _13401_/Y sky130_fd_sc_hd__nand2_1
X_10613_ _19058_/Q _19026_/Q _10613_/S vssd1 vssd1 vccd1 vccd1 _10613_/X sky130_fd_sc_hd__mux2_1
X_14381_ _18233_/Q _16522_/A0 _14382_/S vssd1 vssd1 vccd1 vccd1 _18233_/D sky130_fd_sc_hd__mux2_1
X_11593_ _19066_/Q _19034_/Q _11613_/S vssd1 vssd1 vccd1 vccd1 _11593_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16120_ _16140_/A1 _16119_/Y _16128_/B1 vssd1 vssd1 vccd1 vccd1 _18762_/D sky130_fd_sc_hd__a21oi_1
X_13332_ _17932_/Q _13742_/A2 _13331_/X _14029_/C1 vssd1 vssd1 vccd1 vccd1 _17932_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10544_ _18867_/Q _10613_/S vssd1 vssd1 vccd1 vccd1 _10544_/X sky130_fd_sc_hd__or2_1
XFILLER_259_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16051_ _18730_/Q _18737_/Q _16051_/S vssd1 vssd1 vccd1 vccd1 _16052_/B sky130_fd_sc_hd__mux2_1
X_13263_ _13263_/A _13263_/B vssd1 vssd1 vccd1 vccd1 _13263_/Y sky130_fd_sc_hd__nor2_1
X_10475_ _10850_/A1 _19579_/Q _10840_/S _19611_/Q vssd1 vssd1 vccd1 vccd1 _10475_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15002_ _17821_/Q _15002_/B vssd1 vssd1 vccd1 vccd1 _15002_/X sky130_fd_sc_hd__or2_1
X_12214_ _17869_/Q _12216_/C _12213_/Y vssd1 vssd1 vccd1 vccd1 _17869_/D sky130_fd_sc_hd__o21a_1
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13194_ _13093_/Y _13193_/Y _13194_/S vssd1 vssd1 vccd1 vccd1 _13194_/X sky130_fd_sc_hd__mux2_2
XFILLER_108_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12145_ _17330_/A _12145_/B _12146_/B vssd1 vssd1 vccd1 vccd1 _17843_/D sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19148_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_111_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16953_ _18769_/Q _16965_/A2 _16965_/B1 input234/X _16965_/C1 vssd1 vssd1 vccd1 vccd1
+ _16953_/X sky130_fd_sc_hd__a221o_1
XFILLER_150_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12076_ _17913_/Q _12086_/A2 _12075_/X _17419_/C1 vssd1 vssd1 vccd1 vccd1 _17815_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15904_ _18677_/Q _15910_/A2 _15903_/X _15904_/C1 vssd1 vssd1 vccd1 vccd1 _18677_/D
+ sky130_fd_sc_hd__o211a_1
X_11027_ _18254_/Q _18829_/Q _18457_/Q _18358_/Q _11513_/B2 _11510_/S1 vssd1 vssd1
+ vccd1 vccd1 _11028_/B sky130_fd_sc_hd__mux4_1
X_16884_ _16972_/A _16884_/B vssd1 vssd1 vccd1 vccd1 _19305_/D sky130_fd_sc_hd__and2_1
XFILLER_265_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_202_wb_clk_i _19652_/A vssd1 vssd1 vccd1 vccd1 _19216_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18623_ _19225_/CLK _18623_/D vssd1 vssd1 vccd1 vccd1 _18623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _15835_/A _15835_/B _15835_/C vssd1 vssd1 vccd1 vccd1 _15835_/X sky130_fd_sc_hd__and3_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18554_ _19146_/CLK _18554_/D vssd1 vssd1 vccd1 vccd1 _18554_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _15766_/A _15766_/B vssd1 vssd1 vccd1 vccd1 _15770_/A sky130_fd_sc_hd__and2_1
X_12978_ _13303_/B2 _12963_/X _12966_/X _12977_/X vssd1 vssd1 vccd1 vccd1 _12978_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_45_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _11668_/Y _17520_/A2 _17532_/A2 _17813_/Q _17538_/A vssd1 vssd1 vccd1 vccd1
+ _17505_/X sky130_fd_sc_hd__a221o_1
XFILLER_233_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14717_ input65/X input70/X _14784_/S vssd1 vssd1 vccd1 vccd1 _14718_/B sky130_fd_sc_hd__mux2_8
X_18485_ _19323_/CLK _18485_/D vssd1 vssd1 vccd1 vccd1 _18485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11929_ _11810_/A _11944_/A1 _11810_/C _11959_/A2 input246/X vssd1 vssd1 vccd1 vccd1
+ _11929_/X sky130_fd_sc_hd__a32o_4
XFILLER_233_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15697_ _19482_/Q _15696_/Y _15716_/S vssd1 vssd1 vccd1 vccd1 _15697_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_470 _18380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_481 input233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17436_ _18571_/Q _17527_/A1 _17546_/A2 vssd1 vssd1 vccd1 vccd1 _17436_/X sky130_fd_sc_hd__o21a_1
XANTENNA_492 _18120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14648_ _17707_/A0 _18454_/Q _14648_/S vssd1 vssd1 vccd1 vccd1 _18454_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_17 _14919_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_28 _17181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17367_ _19481_/Q _17196_/B _17379_/S vssd1 vssd1 vccd1 vccd1 _17368_/B sky130_fd_sc_hd__mux2_1
XANTENNA_39 _09139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14579_ _18398_/Q _14589_/A2 _14589_/B1 input27/X vssd1 vssd1 vccd1 vccd1 _14580_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19106_ _19138_/CLK _19106_/D vssd1 vssd1 vccd1 vccd1 _19106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16318_ _17716_/A0 _18931_/Q _16320_/S vssd1 vssd1 vccd1 vccd1 _18931_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17298_ _19450_/Q _17307_/B vssd1 vssd1 vccd1 vccd1 _17298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19037_ _19133_/CLK _19037_/D vssd1 vssd1 vccd1 vccd1 _19037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16249_ _16580_/A0 _18864_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _18864_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09623_ _11161_/S _09622_/X _09106_/B vssd1 vssd1 vccd1 vccd1 _09623_/X sky130_fd_sc_hd__o21a_1
XFILLER_256_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09554_ _09553_/A _09547_/Y _09553_/Y _09350_/S vssd1 vssd1 vccd1 vccd1 _09554_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_243_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09485_ _09908_/A1 _09232_/A _09484_/X _09656_/B1 _18403_/Q vssd1 vssd1 vccd1 vccd1
+ _10084_/B sky130_fd_sc_hd__o32a_1
XFILLER_197_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_77_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19208_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_169_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _10315_/S _10259_/X _10260_/B1 vssd1 vssd1 vccd1 vccd1 _10260_/X sky130_fd_sc_hd__o21a_1
XFILLER_164_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10191_ _18655_/Q _18077_/Q _19096_/Q _19000_/Q _10090_/S _11001_/C1 vssd1 vssd1
+ vccd1 vccd1 _10191_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1305 _12272_/X vssd1 vssd1 vccd1 vccd1 _12276_/A sky130_fd_sc_hd__buf_6
Xfanout1316 _12417_/B1 vssd1 vssd1 vccd1 vccd1 _12429_/B1 sky130_fd_sc_hd__buf_6
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1327 _09098_/Y vssd1 vssd1 vccd1 vccd1 _10260_/B1 sky130_fd_sc_hd__clkbuf_16
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1338 _11459_/A1 vssd1 vssd1 vccd1 vccd1 _10409_/A sky130_fd_sc_hd__buf_8
XFILLER_120_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1349 _09919_/C1 vssd1 vssd1 vccd1 vccd1 _09845_/S sky130_fd_sc_hd__buf_8
X_13950_ _19359_/Q _13950_/A2 _13950_/B1 _19487_/Q _13950_/C1 vssd1 vssd1 vccd1 vccd1
+ _13950_/X sky130_fd_sc_hd__a221o_1
XFILLER_275_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12901_ _13312_/A _14141_/C vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__and2_1
XFILLER_19_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13881_ _19421_/Q _13948_/A2 _13948_/B1 vssd1 vssd1 vccd1 vccd1 _13881_/X sky130_fd_sc_hd__a21o_1
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15620_ _15620_/A _15620_/B _15638_/D vssd1 vssd1 vccd1 vccd1 _15620_/X sky130_fd_sc_hd__or3_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _13314_/S _12831_/Y _12745_/X vssd1 vssd1 vccd1 vccd1 _12833_/A sky130_fd_sc_hd__a21boi_1
XFILLER_74_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _18121_/Q _15763_/A2 _15550_/X _13899_/A vssd1 vssd1 vccd1 vccd1 _15553_/B
+ sky130_fd_sc_hd__a2bb2o_4
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12763_ _13237_/B1 _15216_/A1 _15259_/B _18101_/Q vssd1 vssd1 vccd1 vccd1 _12763_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_243_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _17704_/A0 _18352_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _18352_/D sky130_fd_sc_hd__mux2_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _18524_/Q _18525_/Q _18526_/Q _18527_/Q vssd1 vssd1 vccd1 vccd1 _11715_/D
+ sky130_fd_sc_hd__or4_4
X_18270_ _18272_/CLK _18270_/D vssd1 vssd1 vccd1 vccd1 _18270_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _15484_/A _15484_/C _15484_/B vssd1 vssd1 vccd1 vccd1 _15482_/Y sky130_fd_sc_hd__a21oi_2
X_12694_ _12612_/B _12650_/B _12729_/B vssd1 vssd1 vccd1 vccd1 _12694_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _18101_/Q _17389_/B1 _17394_/A _17256_/B vssd1 vssd1 vccd1 vccd1 _17221_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14433_ _18572_/Q _16052_/A vssd1 vssd1 vccd1 vccd1 _18285_/D sky130_fd_sc_hd__and2_1
XFILLER_230_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11645_ _11728_/A _13904_/B _17531_/A _11645_/D vssd1 vssd1 vccd1 vccd1 _11666_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_230_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17152_ _19402_/Q _17124_/B _17443_/A _17158_/B2 vssd1 vssd1 vccd1 vccd1 _17153_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14364_ _18216_/Q _17671_/A0 _14382_/S vssd1 vssd1 vccd1 vccd1 _18216_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 core_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
X_11576_ _18625_/Q _18196_/Q _11576_/S vssd1 vssd1 vccd1 vccd1 _11576_/X sky130_fd_sc_hd__mux2_1
Xinput26 core_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput37 core_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_2
X_16103_ _18754_/Q _16141_/B vssd1 vssd1 vccd1 vccd1 _16103_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput48 dout0[14] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
X_13315_ _12952_/Y _13314_/X _13315_/S vssd1 vssd1 vccd1 vccd1 _13315_/X sky130_fd_sc_hd__mux2_4
Xinput59 dout0[24] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10527_ _10527_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _11545_/B sky130_fd_sc_hd__and2_2
X_17083_ _19375_/Q _17107_/B vssd1 vssd1 vccd1 vccd1 _17083_/X sky130_fd_sc_hd__or2_1
XFILLER_155_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14295_ _17713_/A0 _18154_/Q _14305_/S vssd1 vssd1 vccd1 vccd1 _18154_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16034_ _18737_/Q _18729_/Q _16034_/S vssd1 vssd1 vccd1 vccd1 _16034_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10458_ _10456_/X _10457_/X _08946_/B vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__a21o_1
X_13246_ _19338_/Q _13246_/A2 _13246_/B1 _19466_/Q _12570_/C vssd1 vssd1 vccd1 vccd1
+ _13246_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13177_ _17863_/Q _13945_/A2 _13166_/X _13945_/B2 _13952_/B1 vssd1 vssd1 vccd1 vccd1
+ _13177_/X sky130_fd_sc_hd__a221o_1
X_10389_ _19061_/Q _19029_/Q _10467_/S vssd1 vssd1 vccd1 vccd1 _10389_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12128_ _17836_/Q _17837_/Q _12128_/C vssd1 vssd1 vccd1 vccd1 _12130_/B sky130_fd_sc_hd__and3_1
X_17985_ _19587_/CLK _17985_/D vssd1 vssd1 vccd1 vccd1 _17985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1850 _16904_/A vssd1 vssd1 vccd1 vccd1 _16968_/A sky130_fd_sc_hd__buf_4
X_16936_ _17342_/A _16936_/B vssd1 vssd1 vccd1 vccd1 _19318_/D sky130_fd_sc_hd__and2_1
X_12059_ _17807_/Q _12073_/B vssd1 vssd1 vccd1 vccd1 _12059_/X sky130_fd_sc_hd__or2_1
Xfanout1861 _15910_/C1 vssd1 vssd1 vccd1 vccd1 _15904_/C1 sky130_fd_sc_hd__buf_4
XFILLER_270_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1872 _17285_/A vssd1 vssd1 vccd1 vccd1 _17198_/A sky130_fd_sc_hd__buf_4
Xfanout1883 fanout1905/X vssd1 vssd1 vccd1 vccd1 _12243_/A sky130_fd_sc_hd__buf_4
XFILLER_37_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1894 _16803_/A vssd1 vssd1 vccd1 vccd1 _16808_/A sky130_fd_sc_hd__buf_4
XFILLER_38_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16867_ _16892_/A _16867_/B vssd1 vssd1 vccd1 vccd1 _19301_/D sky130_fd_sc_hd__and2_1
XFILLER_93_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18606_ _19630_/CLK _18606_/D vssd1 vssd1 vccd1 vccd1 _18606_/Q sky130_fd_sc_hd__dfxtp_1
X_15818_ _18610_/Q _16542_/A0 _15829_/S vssd1 vssd1 vccd1 vccd1 _18610_/D sky130_fd_sc_hd__mux2_1
XFILLER_93_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19586_ _19586_/CLK _19586_/D vssd1 vssd1 vccd1 vccd1 _19586_/Q sky130_fd_sc_hd__dfxtp_1
X_16798_ _19287_/Q _16799_/C _19288_/Q vssd1 vssd1 vccd1 vccd1 _16800_/B sky130_fd_sc_hd__a21oi_1
XFILLER_92_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18537_ _19591_/CLK _18537_/D vssd1 vssd1 vccd1 vccd1 _18537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15749_ _15749_/A _15749_/B vssd1 vssd1 vccd1 vccd1 _15749_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_33_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09270_ _09136_/S _09269_/X _09268_/X _09914_/C1 vssd1 vssd1 vccd1 vccd1 _09274_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18468_ _19647_/CLK _18468_/D vssd1 vssd1 vccd1 vccd1 _18468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17419_ _19495_/Q _17453_/B _17417_/X _17418_/Y _17419_/C1 vssd1 vssd1 vccd1 vccd1
+ _19495_/D sky130_fd_sc_hd__o221a_1
XFILLER_166_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18399_ _19466_/CLK _18399_/D vssd1 vssd1 vccd1 vccd1 _18399_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_147_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_195_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19219_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_124_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18517_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08985_ _11053_/A _08964_/Y _08970_/Y _08977_/Y _08984_/X vssd1 vssd1 vccd1 vccd1
+ _08985_/X sky130_fd_sc_hd__o32a_4
XFILLER_87_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09606_ _11199_/S1 _09595_/X _09605_/X _11516_/B1 vssd1 vssd1 vccd1 vccd1 _09606_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09537_ _09845_/S _09536_/X _09106_/B vssd1 vssd1 vccd1 vccd1 _09537_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09468_ _09441_/X _09444_/X _10180_/A vssd1 vssd1 vccd1 vccd1 _09468_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09399_ _11518_/B2 _09334_/X _09398_/X _09523_/A vssd1 vssd1 vccd1 vccd1 _15259_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11430_ _11511_/A _11429_/X _11495_/B1 vssd1 vssd1 vccd1 vccd1 _11431_/B sky130_fd_sc_hd__a21o_1
XFILLER_177_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11361_ _11359_/X _11360_/X _11361_/S vssd1 vssd1 vccd1 vccd1 _11361_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10312_ _17947_/Q _08946_/Y _10311_/X _11451_/B2 vssd1 vssd1 vccd1 vccd1 _10312_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_138_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13100_ _13100_/A _13100_/B vssd1 vssd1 vccd1 vccd1 _17926_/D sky130_fd_sc_hd__and2_1
XFILLER_180_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14080_ _17696_/A0 _18020_/Q _14104_/S vssd1 vssd1 vccd1 vccd1 _18020_/D sky130_fd_sc_hd__mux2_1
X_11292_ _11292_/A _12595_/B vssd1 vssd1 vccd1 vccd1 _11293_/B sky130_fd_sc_hd__and2_2
XFILLER_106_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10243_ _10243_/A _10243_/B vssd1 vssd1 vccd1 vccd1 _10243_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13031_ _13254_/B2 _11740_/Y _12761_/B _13030_/Y _09866_/B vssd1 vssd1 vccd1 vccd1
+ _13051_/B sky130_fd_sc_hd__a221o_1
XFILLER_191_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10174_ _18623_/Q _18194_/Q _10176_/S vssd1 vssd1 vccd1 vccd1 _10174_/X sky130_fd_sc_hd__mux2_1
Xfanout1102 _15102_/Y vssd1 vssd1 vccd1 vccd1 _17556_/A sky130_fd_sc_hd__buf_6
XFILLER_279_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1113 _12454_/X vssd1 vssd1 vccd1 vccd1 _13637_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1124 _12436_/X vssd1 vssd1 vccd1 vccd1 _13791_/A sky130_fd_sc_hd__buf_4
XFILLER_121_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1135 _12319_/Y vssd1 vssd1 vccd1 vccd1 _13970_/B2 sky130_fd_sc_hd__buf_4
XFILLER_120_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17770_ _19612_/CLK _17770_/D vssd1 vssd1 vccd1 vccd1 _17770_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1146 _10194_/C1 vssd1 vssd1 vccd1 vccd1 _09611_/A sky130_fd_sc_hd__buf_12
XFILLER_78_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1157 _16002_/C1 vssd1 vssd1 vccd1 vccd1 _16004_/C1 sky130_fd_sc_hd__clkbuf_8
X_14982_ _17819_/Q _14982_/B vssd1 vssd1 vccd1 vccd1 _14982_/X sky130_fd_sc_hd__or2_1
Xfanout1168 _15851_/Y vssd1 vssd1 vccd1 vccd1 _15903_/B1 sky130_fd_sc_hd__buf_2
XFILLER_248_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1179 _15502_/B vssd1 vssd1 vccd1 vccd1 _15111_/A sky130_fd_sc_hd__buf_4
X_16721_ _19259_/Q _16723_/C _19260_/Q vssd1 vssd1 vccd1 vccd1 _16724_/B sky130_fd_sc_hd__a21oi_1
XFILLER_75_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13933_ _18131_/Q _13934_/B vssd1 vssd1 vccd1 vccd1 _13969_/B sky130_fd_sc_hd__nand2_2
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19440_ _19506_/CLK _19440_/D vssd1 vssd1 vccd1 vccd1 _19440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16652_ _19240_/Q _19239_/Q _19236_/Q _19235_/Q vssd1 vssd1 vccd1 vccd1 _16653_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13864_ _13860_/A _12837_/B _13862_/Y _13863_/X vssd1 vssd1 vccd1 vccd1 _13864_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15603_ _18584_/Q _15621_/C vssd1 vssd1 vccd1 vccd1 _15603_/Y sky130_fd_sc_hd__nand2_1
X_19371_ _19502_/CLK _19371_/D vssd1 vssd1 vccd1 vccd1 _19371_/Q sky130_fd_sc_hd__dfxtp_1
X_12815_ _12815_/A vssd1 vssd1 vccd1 vccd1 _12815_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16583_ _17683_/A0 _19187_/Q _16585_/S vssd1 vssd1 vccd1 vccd1 _19187_/D sky130_fd_sc_hd__mux2_1
X_13795_ _13761_/B _14151_/B _13892_/B1 vssd1 vssd1 vccd1 vccd1 _13795_/X sky130_fd_sc_hd__a21o_1
X_18322_ _19146_/CLK _18322_/D vssd1 vssd1 vccd1 vccd1 _18322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _18581_/Q _15561_/C _15537_/B1 vssd1 vssd1 vccd1 vccd1 _15535_/B sky130_fd_sc_hd__o21ai_1
XFILLER_188_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12746_ _13134_/S _12746_/B vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__or2_2
XFILLER_203_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _18613_/CLK _18253_/D vssd1 vssd1 vccd1 vccd1 _18253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15465_ _18578_/Q _18577_/Q _15465_/C vssd1 vssd1 vccd1 vccd1 _15512_/C sky130_fd_sc_hd__and3_2
X_12677_ _11212_/Y _12595_/B _12733_/S vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17204_ _17210_/A _17204_/B vssd1 vssd1 vccd1 vccd1 _19419_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14416_ _16292_/A0 _18267_/Q _14416_/S vssd1 vssd1 vccd1 vccd1 _18267_/D sky130_fd_sc_hd__mux2_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18184_ _18613_/CLK _18184_/D vssd1 vssd1 vccd1 vccd1 _18184_/Q sky130_fd_sc_hd__dfxtp_1
X_11628_ _11628_/A _13962_/A vssd1 vssd1 vccd1 vccd1 _11629_/B sky130_fd_sc_hd__nand2_2
XFILLER_191_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15396_ _19469_/Q _19403_/Q vssd1 vssd1 vccd1 vccd1 _15398_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17135_ _17141_/A _17135_/B vssd1 vssd1 vccd1 vccd1 _19396_/D sky130_fd_sc_hd__nor2_1
X_14347_ _14423_/B _14347_/B vssd1 vssd1 vccd1 vccd1 _18202_/D sky130_fd_sc_hd__nor2_4
X_11559_ _18563_/Q _18438_/Q _18047_/Q _18015_/Q _11581_/S _11559_/S1 vssd1 vssd1
+ vccd1 vccd1 _11559_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17066_ _17571_/A _17074_/A2 _17065_/X _17346_/A vssd1 vssd1 vccd1 vccd1 _19366_/D
+ sky130_fd_sc_hd__o211a_1
X_14278_ _16431_/A1 _18137_/Q _14304_/S vssd1 vssd1 vccd1 vccd1 _18137_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16017_ _18724_/Q _16019_/A2 _16016_/X _14197_/A vssd1 vssd1 vccd1 vccd1 _18724_/D
+ sky130_fd_sc_hd__o211a_1
X_13229_ _13047_/Y _13228_/X _13390_/S vssd1 vssd1 vccd1 vccd1 _13229_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_6__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_6__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_97_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17968_ _18627_/CLK _17968_/D vssd1 vssd1 vccd1 vccd1 _17968_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1680 _09854_/A vssd1 vssd1 vccd1 vccd1 _11565_/A1 sky130_fd_sc_hd__buf_6
XFILLER_214_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16919_ _19314_/Q _17175_/B _16927_/S vssd1 vssd1 vccd1 vccd1 _16920_/B sky130_fd_sc_hd__mux2_1
Xfanout1691 _11404_/A1 vssd1 vssd1 vccd1 vccd1 _11017_/A1 sky130_fd_sc_hd__buf_6
XFILLER_77_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17899_ _18881_/CLK _17899_/D vssd1 vssd1 vccd1 vccd1 _17899_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_254_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19638_ _19638_/CLK _19638_/D vssd1 vssd1 vccd1 vccd1 _19638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19569_ _19601_/CLK _19569_/D vssd1 vssd1 vccd1 vccd1 _19569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09322_ _11218_/A _09986_/C vssd1 vssd1 vccd1 vccd1 _09322_/X sky130_fd_sc_hd__or2_1
XFILLER_34_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09253_ _09272_/A1 _17767_/Q _09269_/S _18316_/Q _09135_/S vssd1 vssd1 vccd1 vccd1
+ _09253_/X sky130_fd_sc_hd__o221a_1
XFILLER_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09184_ _11389_/A1 _19141_/Q _09181_/S _19109_/Q _10335_/S vssd1 vssd1 vccd1 vccd1
+ _09184_/X sky130_fd_sc_hd__o221a_1
XFILLER_175_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput205 localMemory_wb_adr_i[23] vssd1 vssd1 vccd1 vccd1 input205/X sky130_fd_sc_hd__clkbuf_8
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput216 localMemory_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input216/X sky130_fd_sc_hd__buf_8
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput227 localMemory_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input227/X sky130_fd_sc_hd__clkbuf_16
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput238 localMemory_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 input238/X sky130_fd_sc_hd__buf_12
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ _18854_/Q _18886_/Q _19046_/Q _19014_/Q _08968_/S0 _09978_/A1 vssd1 vssd1
+ vccd1 vccd1 _08968_/X sky130_fd_sc_hd__mux4_1
Xinput249 localMemory_wb_sel_i[2] vssd1 vssd1 vccd1 vccd1 input249/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08899_ _08899_/A _12023_/A vssd1 vssd1 vccd1 vccd1 _08899_/Y sky130_fd_sc_hd__nor2_8
XFILLER_217_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10930_ _10928_/X _10929_/X _10930_/S vssd1 vssd1 vccd1 vccd1 _10930_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_92_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18776_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10861_ _18256_/Q _10853_/S _10785_/A _10860_/X vssd1 vssd1 vccd1 vccd1 _10861_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_21_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18875_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_204_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12600_/A _12600_/B vssd1 vssd1 vccd1 vccd1 _13225_/B sky130_fd_sc_hd__and2_1
XFILLER_25_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _17939_/Q _13742_/A2 _13579_/X _14177_/A vssd1 vssd1 vccd1 vccd1 _17939_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10792_ _10532_/A _10792_/A2 _10791_/X vssd1 vssd1 vccd1 vccd1 _11860_/A sky130_fd_sc_hd__o21ai_1
XFILLER_231_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12531_ _19360_/Q _13925_/S _12527_/X _12530_/X vssd1 vssd1 vccd1 vccd1 _12531_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15250_ _15416_/A _15250_/B _15250_/C vssd1 vssd1 vccd1 vccd1 _15250_/X sky130_fd_sc_hd__or3_1
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12462_ _16821_/A _14004_/A _14992_/A1 vssd1 vssd1 vccd1 vccd1 _12577_/A sky130_fd_sc_hd__a21oi_4
XFILLER_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14201_ _14203_/A _14201_/B vssd1 vssd1 vccd1 vccd1 _18098_/D sky130_fd_sc_hd__and2_1
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11413_ _18545_/Q _18420_/Q _18029_/Q _17997_/Q _11426_/B2 _11510_/S1 vssd1 vssd1
+ vccd1 vccd1 _11413_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15181_ _18566_/Q _18565_/Q _18564_/Q vssd1 vssd1 vccd1 vccd1 _15224_/C sky130_fd_sc_hd__and3_2
X_12393_ _12429_/A1 _09236_/A _09149_/X _12417_/B1 _18391_/Q vssd1 vssd1 vccd1 vccd1
+ _12394_/B sky130_fd_sc_hd__o32ai_4
XFILLER_165_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14132_ _16549_/A0 _18071_/Q _14140_/S vssd1 vssd1 vccd1 vccd1 _18071_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11344_ _11360_/A1 _19209_/Q _19177_/Q _11360_/B2 vssd1 vssd1 vccd1 vccd1 _11344_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18940_ _19201_/CLK _18940_/D vssd1 vssd1 vccd1 vccd1 _18940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14063_ _17680_/A0 _18005_/Q _14073_/S vssd1 vssd1 vccd1 vccd1 _18005_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11275_ _11282_/A _11275_/B vssd1 vssd1 vccd1 vccd1 _11280_/A sky130_fd_sc_hd__and2_1
XFILLER_267_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13014_ _19527_/Q _13372_/S vssd1 vssd1 vccd1 vccd1 _13014_/X sky130_fd_sc_hd__or2_1
X_10226_ _10222_/X _10225_/X _10301_/S vssd1 vssd1 vccd1 vccd1 _10226_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18871_ _19614_/CLK _18871_/D vssd1 vssd1 vccd1 vccd1 _18871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17822_ _18201_/CLK _17822_/D vssd1 vssd1 vccd1 vccd1 _17822_/Q sky130_fd_sc_hd__dfxtp_1
X_10157_ _18131_/Q _10156_/Y _13545_/A vssd1 vssd1 vccd1 vccd1 _12660_/B sky130_fd_sc_hd__mux2_4
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17753_ _18653_/Q vssd1 vssd1 vccd1 vccd1 _18653_/D sky130_fd_sc_hd__clkbuf_2
X_10088_ _17950_/Q _08946_/Y _10087_/X _11451_/B2 vssd1 vssd1 vccd1 vccd1 _10089_/B
+ sky130_fd_sc_hd__o22a_4
X_14965_ _18128_/Q _14671_/X _14934_/X _14964_/X vssd1 vssd1 vccd1 vccd1 _14965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16704_ _19254_/Q _19253_/Q _16704_/C vssd1 vssd1 vccd1 vccd1 _16706_/B sky130_fd_sc_hd__and3_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13916_ _13916_/A _13938_/B vssd1 vssd1 vccd1 vccd1 _13916_/X sky130_fd_sc_hd__or2_1
X_17684_ _17684_/A0 _19611_/Q _17690_/S vssd1 vssd1 vccd1 vccd1 _19611_/D sky130_fd_sc_hd__mux2_1
X_14896_ input55/X input90/X _14947_/S vssd1 vssd1 vccd1 vccd1 _14897_/A sky130_fd_sc_hd__mux2_2
XFILLER_74_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16635_ _19234_/Q _16677_/A _16752_/A vssd1 vssd1 vccd1 vccd1 _16635_/Y sky130_fd_sc_hd__a21oi_1
X_19423_ _19519_/CLK _19423_/D vssd1 vssd1 vccd1 vccd1 _19423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13847_ _17883_/Q _13847_/A2 _13845_/X _13928_/A1 vssd1 vssd1 vccd1 vccd1 _13847_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16566_ _17699_/A0 _19170_/Q _16589_/S vssd1 vssd1 vccd1 vccd1 _19170_/D sky130_fd_sc_hd__mux2_1
X_19354_ _19481_/CLK _19354_/D vssd1 vssd1 vccd1 vccd1 _19354_/Q sky130_fd_sc_hd__dfxtp_1
X_13778_ _17849_/Q _13821_/B vssd1 vssd1 vccd1 vccd1 _13778_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18305_ _18593_/CLK _18305_/D vssd1 vssd1 vccd1 vccd1 _18305_/Q sky130_fd_sc_hd__dfxtp_1
X_15517_ _19442_/Q _15661_/B _17214_/A vssd1 vssd1 vccd1 vccd1 _15517_/X sky130_fd_sc_hd__o21a_1
X_19285_ _19285_/CLK _19285_/D vssd1 vssd1 vccd1 vccd1 _19285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12729_ _12729_/A _12729_/B vssd1 vssd1 vccd1 vccd1 _12729_/X sky130_fd_sc_hd__or2_1
X_16497_ _16530_/A0 _19103_/Q _16521_/S vssd1 vssd1 vccd1 vccd1 _19103_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18236_ _18875_/CLK _18236_/D vssd1 vssd1 vccd1 vccd1 _18236_/Q sky130_fd_sc_hd__dfxtp_1
X_15448_ _15447_/B _15439_/X _15446_/X _15447_/Y _17261_/A vssd1 vssd1 vccd1 vccd1
+ _18577_/D sky130_fd_sc_hd__a311oi_1
XFILLER_157_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18167_ _19620_/CLK _18167_/D vssd1 vssd1 vccd1 vccd1 _18167_/Q sky130_fd_sc_hd__dfxtp_1
X_15379_ _18574_/Q _15447_/B _15370_/X _15378_/X _17469_/C1 vssd1 vssd1 vccd1 vccd1
+ _18574_/D sky130_fd_sc_hd__o221a_1
XFILLER_144_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17118_ _17217_/B _17118_/B _16973_/B vssd1 vssd1 vccd1 vccd1 _17118_/X sky130_fd_sc_hd__or3b_2
X_18098_ _18713_/CLK _18098_/D vssd1 vssd1 vccd1 vccd1 _18098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09940_ _10260_/B1 _09931_/X _09935_/X _09939_/X vssd1 vssd1 vccd1 vccd1 _09940_/X
+ sky130_fd_sc_hd__a31o_1
X_17049_ _17381_/C _17591_/D vssd1 vssd1 vccd1 vccd1 _17073_/B sky130_fd_sc_hd__nor2_8
XFILLER_104_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout906 _16458_/S vssd1 vssd1 vccd1 vccd1 _16454_/S sky130_fd_sc_hd__buf_12
Xfanout917 _16288_/S vssd1 vssd1 vccd1 vccd1 _16291_/S sky130_fd_sc_hd__buf_12
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _12766_/A0 _09867_/X _09870_/X vssd1 vssd1 vccd1 vccd1 _09877_/A sky130_fd_sc_hd__a21oi_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout928 _17543_/B1 vssd1 vssd1 vccd1 vccd1 _17532_/A2 sky130_fd_sc_hd__buf_4
XFILLER_225_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout939 _14973_/C1 vssd1 vssd1 vccd1 vccd1 _15003_/C1 sky130_fd_sc_hd__buf_4
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _18778_/Q vssd1 vssd1 vccd1 vccd1 _14424_/A sky130_fd_sc_hd__inv_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09305_ _09303_/X _09304_/X _09374_/S vssd1 vssd1 vccd1 vccd1 _09305_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09236_ _09236_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _09236_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09167_ _19205_/Q _19173_/Q _09344_/S vssd1 vssd1 vccd1 vccd1 _09167_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09098_ _09750_/S _12023_/A vssd1 vssd1 vccd1 vccd1 _09098_/Y sky130_fd_sc_hd__nor2_8
XFILLER_253_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11060_ _13535_/S vssd1 vssd1 vccd1 vccd1 _11060_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_150_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10011_ _18236_/Q _18811_/Q _10840_/S vssd1 vssd1 vccd1 vccd1 _10011_/X sky130_fd_sc_hd__mux2_1
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _17796_/Q _14982_/B vssd1 vssd1 vccd1 vccd1 _14750_/X sky130_fd_sc_hd__or2_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11962_ _18508_/Q _11720_/X _11912_/X _11968_/B2 vssd1 vssd1 vccd1 vccd1 _11962_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _13896_/B2 _13156_/Y _13700_/X vssd1 vssd1 vccd1 vccd1 _13701_/X sky130_fd_sc_hd__o21a_1
XFILLER_260_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10913_ _17939_/Q _08948_/B _10912_/Y _08947_/B vssd1 vssd1 vccd1 vccd1 _10913_/X
+ sky130_fd_sc_hd__o22a_4
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _12292_/C _14681_/B _14681_/C vssd1 vssd1 vccd1 vccd1 _14683_/A sky130_fd_sc_hd__and3b_1
XFILLER_45_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _11820_/Y _11875_/Y _11892_/X vssd1 vssd1 vccd1 vccd1 _11894_/C sky130_fd_sc_hd__o21ai_2
XFILLER_72_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16420_ _16618_/A0 _19029_/Q _16420_/S vssd1 vssd1 vccd1 vccd1 _19029_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13632_ _19349_/Q _13950_/A2 _13950_/B1 _19477_/Q _13950_/C1 vssd1 vssd1 vccd1 vccd1
+ _13632_/X sky130_fd_sc_hd__a221o_1
X_10844_ _11568_/A _10842_/X _10843_/X _11570_/B1 vssd1 vssd1 vccd1 vccd1 _10844_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_25_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16351_ _18963_/Q _10532_/B _16358_/S vssd1 vssd1 vccd1 vccd1 _18963_/D sky130_fd_sc_hd__mux2_1
XFILLER_241_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13563_ _13438_/A _13548_/X _13563_/B1 vssd1 vssd1 vccd1 vccd1 _13563_/X sky130_fd_sc_hd__a21o_1
X_10775_ _11328_/S _10770_/X _10774_/X _11588_/B1 vssd1 vssd1 vccd1 vccd1 _10775_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_200_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15302_ _18571_/Q _15351_/A2 _15296_/X _15301_/X _17469_/C1 vssd1 vssd1 vccd1 vccd1
+ _18571_/D sky130_fd_sc_hd__o221a_1
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12514_ _12514_/A _12514_/B vssd1 vssd1 vccd1 vccd1 _12552_/A sky130_fd_sc_hd__nand2_4
X_19070_ _19114_/CLK _19070_/D vssd1 vssd1 vccd1 vccd1 _19070_/Q sky130_fd_sc_hd__dfxtp_1
X_16282_ _16580_/A0 _18896_/Q _16292_/S vssd1 vssd1 vccd1 vccd1 _18896_/D sky130_fd_sc_hd__mux2_1
X_13494_ _17840_/Q _13846_/B _12548_/X vssd1 vssd1 vccd1 vccd1 _13494_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18021_ _18902_/CLK _18021_/D vssd1 vssd1 vccd1 vccd1 _18021_/Q sky130_fd_sc_hd__dfxtp_1
X_15233_ _15233_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15233_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_139_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12445_ _12445_/A _12445_/B vssd1 vssd1 vccd1 vccd1 _12448_/D sky130_fd_sc_hd__nand2_4
XFILLER_126_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15164_ _19459_/Q _19393_/Q vssd1 vssd1 vccd1 vccd1 _15166_/A sky130_fd_sc_hd__and2_1
XFILLER_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12376_ _12408_/B _12376_/B vssd1 vssd1 vccd1 vccd1 _12376_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14115_ _16532_/A0 _18054_/Q _14131_/S vssd1 vssd1 vccd1 vccd1 _18054_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11327_ _11325_/X _11326_/X _11327_/S vssd1 vssd1 vccd1 vccd1 _11327_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15095_ _19382_/Q _15086_/B input183/X _15094_/X vssd1 vssd1 vccd1 vccd1 _15101_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_119_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14046_ _17696_/A0 _17988_/Q _14070_/S vssd1 vssd1 vccd1 vccd1 _17988_/D sky130_fd_sc_hd__mux2_1
X_18923_ _19634_/CLK _18923_/D vssd1 vssd1 vccd1 vccd1 _18923_/Q sky130_fd_sc_hd__dfxtp_1
X_11258_ _11488_/A _11832_/A vssd1 vssd1 vccd1 vccd1 _11258_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10209_ _10200_/S _10202_/X _10201_/X _10356_/C1 vssd1 vssd1 vccd1 vccd1 _10209_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_192_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18854_ _19206_/CLK _18854_/D vssd1 vssd1 vccd1 vccd1 _18854_/Q sky130_fd_sc_hd__dfxtp_1
X_11189_ _11189_/A _11189_/B vssd1 vssd1 vccd1 vccd1 _11194_/A sky130_fd_sc_hd__and2_1
XFILLER_283_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17805_ _17814_/CLK _17805_/D vssd1 vssd1 vccd1 vccd1 _17805_/Q sky130_fd_sc_hd__dfxtp_2
X_15997_ _18714_/Q _16005_/A2 _15996_/X _14205_/A vssd1 vssd1 vccd1 vccd1 _18714_/D
+ sky130_fd_sc_hd__o211a_1
X_18785_ _19624_/CLK _18785_/D vssd1 vssd1 vccd1 vccd1 _18785_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17736_ _18636_/Q vssd1 vssd1 vccd1 vccd1 _18636_/D sky130_fd_sc_hd__clkbuf_2
X_14948_ _14948_/A vssd1 vssd1 vccd1 vccd1 _14948_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_36_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17667_ _17667_/A0 _19594_/Q _17689_/S vssd1 vssd1 vccd1 vccd1 _19594_/D sky130_fd_sc_hd__mux2_1
X_14879_ _14875_/Y _14878_/X _14879_/B1 vssd1 vssd1 vccd1 vccd1 _14879_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19406_ _19537_/CLK _19406_/D vssd1 vssd1 vccd1 vccd1 _19406_/Q sky130_fd_sc_hd__dfxtp_1
X_16618_ _16618_/A0 _19221_/Q _16618_/S vssd1 vssd1 vccd1 vccd1 _19221_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17598_ _19540_/Q _17622_/A2 _17591_/X _17175_/B _17597_/X vssd1 vssd1 vccd1 vccd1
+ _19540_/D sky130_fd_sc_hd__o221a_1
XFILLER_210_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16549_ _16549_/A0 _19154_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _19154_/D sky130_fd_sc_hd__mux2_1
X_19337_ _19465_/CLK _19337_/D vssd1 vssd1 vccd1 vccd1 _19337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19268_ _19268_/CLK _19268_/D vssd1 vssd1 vccd1 vccd1 _19268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09021_ _11217_/C _11556_/C vssd1 vssd1 vccd1 vccd1 _09021_/X sky130_fd_sc_hd__or2_1
XFILLER_148_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18219_ _19146_/CLK _18219_/D vssd1 vssd1 vccd1 vccd1 _18219_/Q sky130_fd_sc_hd__dfxtp_1
X_19199_ _19622_/CLK _19199_/D vssd1 vssd1 vccd1 vccd1 _19199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09923_ _09683_/A _09915_/X _09916_/X _10260_/B1 _09914_/X vssd1 vssd1 vccd1 vccd1
+ _09923_/X sky130_fd_sc_hd__o311a_1
Xfanout703 _12544_/Y vssd1 vssd1 vccd1 vccd1 _13495_/A2 sky130_fd_sc_hd__buf_4
Xfanout714 _12919_/A2 vssd1 vssd1 vccd1 vccd1 _13847_/A2 sky130_fd_sc_hd__buf_4
XFILLER_59_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout725 _12495_/Y vssd1 vssd1 vccd1 vccd1 _13844_/A2 sky130_fd_sc_hd__buf_4
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout736 _17706_/A0 vssd1 vssd1 vccd1 vccd1 _16606_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout747 _13263_/A vssd1 vssd1 vccd1 vccd1 _13314_/S sky130_fd_sc_hd__buf_4
X_09854_ _09854_/A _19556_/Q _15082_/A vssd1 vssd1 vccd1 vccd1 _09854_/X sky130_fd_sc_hd__or3_1
Xfanout758 _09160_/X vssd1 vssd1 vccd1 vccd1 _17702_/A0 sky130_fd_sc_hd__buf_6
XFILLER_112_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout769 _17658_/Y vssd1 vssd1 vccd1 vccd1 _17690_/S sky130_fd_sc_hd__buf_12
XFILLER_252_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ _18597_/Q _18168_/Q _09797_/S vssd1 vssd1 vccd1 vccd1 _09785_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _11732_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_118 _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _11814_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10560_ _10618_/S _10559_/X _11570_/B1 vssd1 vssd1 vccd1 vccd1 _10560_/X sky130_fd_sc_hd__o21a_1
XFILLER_194_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ _10354_/A1 _18214_/Q _10348_/S _18949_/Q _10205_/S vssd1 vssd1 vccd1 vccd1
+ _09219_/X sky130_fd_sc_hd__o221a_1
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10491_ _18332_/Q _17783_/Q _10500_/S vssd1 vssd1 vccd1 vccd1 _10491_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12230_ _17875_/Q _12232_/C _12229_/Y vssd1 vssd1 vccd1 vccd1 _17875_/D sky130_fd_sc_hd__o21a_1
XFILLER_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12161_ _12243_/A _12161_/B _12162_/B vssd1 vssd1 vccd1 vccd1 _17849_/D sky130_fd_sc_hd__nor3_1
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11112_ _11112_/A _11112_/B vssd1 vssd1 vccd1 vccd1 _11117_/A sky130_fd_sc_hd__and2_1
XFILLER_122_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12092_ _17823_/Q _17824_/Q _12107_/A vssd1 vssd1 vccd1 vccd1 _12092_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_268_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15920_ _15920_/A _15947_/S _15923_/C vssd1 vssd1 vccd1 vccd1 _15920_/X sky130_fd_sc_hd__and3_1
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ _18861_/Q _18893_/Q _19053_/Q _19021_/Q _09290_/S _11503_/S1 vssd1 vssd1
+ vccd1 vccd1 _11043_/X sky130_fd_sc_hd__mux4_1
XFILLER_249_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15851_ _15853_/A _15955_/B vssd1 vssd1 vccd1 vccd1 _15851_/Y sky130_fd_sc_hd__nand2_2
XFILLER_249_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _14964_/B1 _14800_/X _14801_/X _14771_/X vssd1 vssd1 vccd1 vccd1 _14802_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15782_ _15782_/A1 _15781_/X _15782_/B1 vssd1 vssd1 vccd1 vccd1 _15782_/X sky130_fd_sc_hd__a21o_1
X_18570_ _19399_/CLK _18570_/D vssd1 vssd1 vccd1 vccd1 _18570_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_224_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12994_ _12994_/A vssd1 vssd1 vccd1 vccd1 _12994_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14733_ _14992_/A1 _12978_/X _14973_/B1 _18630_/Q _14741_/B vssd1 vssd1 vccd1 vccd1
+ _14733_/X sky130_fd_sc_hd__a221o_1
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17521_ _18588_/Q _17544_/A _17520_/X _08883_/A vssd1 vssd1 vccd1 vccd1 _17521_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_205_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ _11959_/B2 _11882_/B _11882_/C _11945_/B1 input232/X vssd1 vssd1 vccd1 vccd1
+ _11945_/X sky130_fd_sc_hd__a32o_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17452_ _18113_/Q _17463_/A2 _17450_/X _17451_/X vssd1 vssd1 vccd1 vccd1 _17452_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14664_ _17723_/A0 _18470_/Q _14664_/S vssd1 vssd1 vccd1 vccd1 _18470_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11876_ _11804_/X _11875_/A _11901_/B _11837_/X vssd1 vssd1 vccd1 vccd1 _11876_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _17668_/A0 _19012_/Q _16424_/S vssd1 vssd1 vccd1 vccd1 _19012_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13615_ _13615_/A _13615_/B vssd1 vssd1 vccd1 vccd1 _13616_/B sky130_fd_sc_hd__nand2_1
X_10827_ _11365_/B2 _10792_/A2 _10826_/Y _11133_/B2 vssd1 vssd1 vccd1 vccd1 _13623_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_17383_ _19231_/Q _12322_/Y _17129_/Y _17382_/B vssd1 vssd1 vccd1 vccd1 _17383_/X
+ sky130_fd_sc_hd__a22o_1
X_14595_ _14593_/X _14594_/X input9/X _11689_/A vssd1 vssd1 vccd1 vccd1 _14596_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16334_ _18946_/Q _09437_/B _16355_/S vssd1 vssd1 vccd1 vccd1 _18946_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19122_ _19154_/CLK _19122_/D vssd1 vssd1 vccd1 vccd1 _19122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13546_ _17906_/Q _13971_/A2 _13544_/Y _13545_/X _13579_/A vssd1 vssd1 vccd1 vccd1
+ _13546_/X sky130_fd_sc_hd__a221o_4
X_10758_ _17973_/Q _16820_/A3 _11216_/B1 vssd1 vssd1 vccd1 vccd1 _10758_/X sky130_fd_sc_hd__a21o_1
XFILLER_201_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19053_ _19213_/CLK _19053_/D vssd1 vssd1 vccd1 vccd1 _19053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16265_ _16431_/A1 _18879_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _18879_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13477_ _10513_/S _12448_/C _13475_/Y _13476_/X _12762_/B vssd1 vssd1 vccd1 vccd1
+ _13477_/X sky130_fd_sc_hd__a221o_4
XFILLER_127_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10689_ _10685_/X _10688_/X _10689_/S vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__mux2_1
X_18004_ _19649_/CLK _18004_/D vssd1 vssd1 vccd1 vccd1 _18004_/Q sky130_fd_sc_hd__dfxtp_1
X_15216_ _15216_/A1 _15285_/A3 _18107_/Q vssd1 vssd1 vccd1 vccd1 _15216_/X sky130_fd_sc_hd__a21o_1
X_12428_ _17917_/Q _12427_/A _12427_/Y _12428_/C1 vssd1 vssd1 vccd1 vccd1 _17917_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16196_ _17693_/A0 _18812_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _18812_/D sky130_fd_sc_hd__mux2_1
Xoutput306 _11754_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[10] sky130_fd_sc_hd__buf_4
XFILLER_127_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput317 _11764_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[20] sky130_fd_sc_hd__buf_4
Xoutput328 _11741_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[5] sky130_fd_sc_hd__buf_4
X_15147_ _17141_/A _15147_/B vssd1 vssd1 vccd1 vccd1 _15147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12359_ _17894_/Q _12421_/A _12358_/Y _14417_/A vssd1 vssd1 vccd1 vccd1 _17894_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput339 _11831_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[14] sky130_fd_sc_hd__buf_4
XFILLER_236_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15078_ _18562_/Q _16490_/A0 _15078_/S vssd1 vssd1 vccd1 vccd1 _18562_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14029_ _17979_/Q _14028_/A _14028_/Y _14029_/C1 vssd1 vssd1 vccd1 vccd1 _17979_/D
+ sky130_fd_sc_hd__o211a_1
X_18906_ _19055_/CLK _18906_/D vssd1 vssd1 vccd1 vccd1 _18906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18837_ _19055_/CLK _18837_/D vssd1 vssd1 vccd1 vccd1 _18837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09570_ _09908_/A1 _09232_/A _09569_/X _09908_/B1 _18402_/Q vssd1 vssd1 vccd1 vccd1
+ _10162_/B sky130_fd_sc_hd__o32a_1
XFILLER_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18768_ _18772_/CLK _18768_/D vssd1 vssd1 vccd1 vccd1 _18768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_255_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17719_ _17719_/A0 _19645_/Q _17719_/S vssd1 vssd1 vccd1 vccd1 _19645_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18699_ _18700_/CLK _18699_/D vssd1 vssd1 vccd1 vccd1 _18699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_149_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19526_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_282_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09004_ input131/X input166/X _09657_/S vssd1 vssd1 vccd1 vccd1 _09004_/X sky130_fd_sc_hd__mux2_8
XFILLER_136_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout500 _11706_/X vssd1 vssd1 vccd1 vccd1 _11968_/B2 sky130_fd_sc_hd__buf_8
XFILLER_278_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1509 fanout1514/X vssd1 vssd1 vccd1 vccd1 _10128_/B sky130_fd_sc_hd__buf_6
Xfanout511 _17499_/A2 vssd1 vssd1 vccd1 vccd1 _17423_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09906_ input118/X input133/X _09990_/S vssd1 vssd1 vccd1 vccd1 _09907_/B sky130_fd_sc_hd__mux2_8
XFILLER_59_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout522 _15127_/Y vssd1 vssd1 vccd1 vccd1 _15718_/A2 sky130_fd_sc_hd__buf_4
Xfanout533 fanout536/X vssd1 vssd1 vccd1 vccd1 fanout533/X sky130_fd_sc_hd__buf_4
XFILLER_132_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout544 _17129_/A vssd1 vssd1 vccd1 vccd1 _17219_/A sky130_fd_sc_hd__buf_4
Xfanout555 _15122_/Y vssd1 vssd1 vccd1 vccd1 _17157_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_258_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout566 _15132_/X vssd1 vssd1 vccd1 vccd1 _15786_/A2 sky130_fd_sc_hd__buf_6
XFILLER_259_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout577 _12379_/A vssd1 vssd1 vccd1 vccd1 _12349_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09837_ _18845_/Q _18877_/Q _11147_/S vssd1 vssd1 vccd1 vccd1 _09837_/X sky130_fd_sc_hd__mux2_1
Xfanout588 _12073_/B vssd1 vssd1 vccd1 vccd1 _12051_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_274_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout599 _14260_/B vssd1 vssd1 vccd1 vccd1 _14266_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09768_ _09768_/A _09768_/B vssd1 vssd1 vccd1 vccd1 _09768_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _09696_/X _09697_/Y _09946_/B1 vssd1 vssd1 vccd1 vccd1 _12609_/A sky130_fd_sc_hd__a21o_2
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _14522_/A2 _15039_/B vssd1 vssd1 vccd1 vccd1 _11730_/Y sky130_fd_sc_hd__nand2b_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _15082_/B _15120_/B vssd1 vssd1 vccd1 vccd1 _11774_/B sky130_fd_sc_hd__and2_4
XFILLER_230_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13400_ _15429_/A2 _13396_/X _13399_/X _13936_/B2 vssd1 vssd1 vccd1 vccd1 _13401_/B
+ sky130_fd_sc_hd__a22o_1
X_10612_ _10610_/X _10611_/X _10633_/A vssd1 vssd1 vccd1 vccd1 _10612_/X sky130_fd_sc_hd__mux2_1
X_14380_ _18232_/Q _16488_/A0 _14380_/S vssd1 vssd1 vccd1 vccd1 _18232_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11592_ _15549_/A _11591_/X _11592_/S vssd1 vssd1 vccd1 vccd1 _11628_/A sky130_fd_sc_hd__mux2_4
XFILLER_211_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _17900_/Q _12448_/C _13329_/Y _13330_/Y _13808_/C1 vssd1 vssd1 vccd1 vccd1
+ _13331_/X sky130_fd_sc_hd__a221o_4
X_10543_ _10541_/X _10542_/X _10618_/S vssd1 vssd1 vccd1 vccd1 _10543_/X sky130_fd_sc_hd__mux2_4
XFILLER_155_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16050_ _16052_/A _16050_/B vssd1 vssd1 vccd1 vccd1 _18736_/D sky130_fd_sc_hd__and2_1
X_13262_ _13312_/A _13261_/X _13909_/B1 _13258_/Y vssd1 vssd1 vccd1 vccd1 _13262_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire989 wire989/A vssd1 vssd1 vccd1 vccd1 wire989/X sky130_fd_sc_hd__buf_6
X_10474_ _18557_/Q _18432_/Q _18041_/Q _18009_/Q _10840_/S _10918_/C1 vssd1 vssd1
+ vccd1 vccd1 _10474_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15001_ _18501_/Q _15001_/A2 _15000_/Y _16787_/A vssd1 vssd1 vccd1 vccd1 _18501_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12213_ _17869_/Q _12216_/C _12219_/A vssd1 vssd1 vccd1 vccd1 _12213_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13193_ _13193_/A vssd1 vssd1 vccd1 vccd1 _13193_/Y sky130_fd_sc_hd__inv_2
XFILLER_269_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12144_ _17842_/Q _17843_/Q _12144_/C vssd1 vssd1 vccd1 vccd1 _12146_/B sky130_fd_sc_hd__and3_1
XFILLER_2_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16952_ _16960_/A _16952_/B vssd1 vssd1 vccd1 vccd1 _19322_/D sky130_fd_sc_hd__and2_1
X_12075_ _17815_/Q _12085_/B vssd1 vssd1 vccd1 vccd1 _12075_/X sky130_fd_sc_hd__or2_1
XFILLER_111_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15903_ _18676_/Q _15906_/A2 _15903_/B1 _15902_/X vssd1 vssd1 vccd1 vccd1 _15903_/X
+ sky130_fd_sc_hd__a211o_1
X_11026_ _17906_/Q _11135_/S _11181_/B1 _11025_/Y vssd1 vssd1 vccd1 vccd1 _12594_/A
+ sky130_fd_sc_hd__o22a_2
X_16883_ _19305_/Q _17577_/A _16971_/S vssd1 vssd1 vccd1 vccd1 _16884_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18622_ _19646_/CLK _18622_/D vssd1 vssd1 vccd1 vccd1 _18622_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _16819_/A _15834_/B _15834_/C vssd1 vssd1 vccd1 vccd1 _15843_/A sky130_fd_sc_hd__nor3_4
XFILLER_265_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18553_ _19600_/CLK _18553_/D vssd1 vssd1 vccd1 vccd1 _18553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12977_ _12977_/A _12977_/B vssd1 vssd1 vccd1 vccd1 _12977_/X sky130_fd_sc_hd__or2_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _15787_/A _15765_/B vssd1 vssd1 vccd1 vccd1 _15766_/B sky130_fd_sc_hd__or2_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17504_ _19512_/Q _17523_/B _17502_/X _17503_/Y _17592_/B vssd1 vssd1 vccd1 vccd1
+ _19512_/D sky130_fd_sc_hd__o221a_1
XFILLER_221_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14716_ _18658_/Q _16819_/B _14685_/X _14875_/A1 _14715_/X vssd1 vssd1 vccd1 vccd1
+ _14716_/X sky130_fd_sc_hd__a311o_1
X_11928_ _11810_/A _11944_/A1 _11806_/C _11959_/A2 input245/X vssd1 vssd1 vccd1 vccd1
+ _11928_/X sky130_fd_sc_hd__a32o_4
X_18484_ _18517_/CLK _18484_/D vssd1 vssd1 vccd1 vccd1 _18484_/Q sky130_fd_sc_hd__dfxtp_1
X_15696_ _15696_/A _15696_/B vssd1 vssd1 vccd1 vccd1 _15696_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_460 _18373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_471 _18731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ _16606_/A0 _18453_/Q _14664_/S vssd1 vssd1 vccd1 vccd1 _18453_/D sky130_fd_sc_hd__mux2_1
XANTENNA_482 input237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17435_ _11751_/Y _17475_/A2 _17475_/B1 _17799_/Q _15116_/B vssd1 vssd1 vccd1 vccd1
+ _17435_/X sky130_fd_sc_hd__a221o_1
XFILLER_205_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_493 _18131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11859_ _11859_/A _11859_/B vssd1 vssd1 vccd1 vccd1 _11875_/A sky130_fd_sc_hd__nand2_8
XFILLER_268_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 _14919_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_29 _17199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17366_ _17366_/A _17366_/B vssd1 vssd1 vccd1 vccd1 _19480_/D sky130_fd_sc_hd__and2_1
X_14578_ _14592_/A _14578_/B vssd1 vssd1 vccd1 vccd1 _18397_/D sky130_fd_sc_hd__or2_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19105_ _19147_/CLK _19105_/D vssd1 vssd1 vccd1 vccd1 _19105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16317_ _17715_/A0 _18930_/Q _16320_/S vssd1 vssd1 vccd1 vccd1 _18930_/D sky130_fd_sc_hd__mux2_1
X_13529_ _13930_/A1 _13515_/Y _13930_/B1 vssd1 vssd1 vccd1 vccd1 _13529_/Y sky130_fd_sc_hd__o21ai_1
X_17297_ _17295_/Y _17296_/X _17198_/A vssd1 vssd1 vccd1 vccd1 _19449_/D sky130_fd_sc_hd__a21oi_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19036_ _19196_/CLK _19036_/D vssd1 vssd1 vccd1 vccd1 _19036_/Q sky130_fd_sc_hd__dfxtp_1
X_16248_ _17712_/A0 _18863_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _18863_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16179_ _17709_/A0 _18796_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _18796_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09622_ _18631_/Q _18053_/Q _19072_/Q _18976_/Q _11171_/S _11156_/C1 vssd1 vssd1
+ vccd1 vccd1 _09622_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09553_ _09553_/A _09553_/B vssd1 vssd1 vccd1 vccd1 _09553_/Y sky130_fd_sc_hd__nor2_1
XFILLER_270_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09484_ input130/X input165/X _09655_/S vssd1 vssd1 vccd1 vccd1 _09484_/X sky130_fd_sc_hd__mux2_8
XFILLER_23_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18880_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10190_ _10336_/A _10190_/B vssd1 vssd1 vccd1 vccd1 _10190_/X sky130_fd_sc_hd__or2_2
XFILLER_274_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1306 _15941_/S vssd1 vssd1 vccd1 vccd1 _15905_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_160_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1317 _12420_/B1 vssd1 vssd1 vccd1 vccd1 _12417_/B1 sky130_fd_sc_hd__buf_8
XFILLER_120_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1328 _10633_/A vssd1 vssd1 vccd1 vccd1 _10785_/A sky130_fd_sc_hd__buf_8
XFILLER_278_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1339 _10004_/A1 vssd1 vssd1 vccd1 vccd1 _11459_/A1 sky130_fd_sc_hd__buf_6
XFILLER_219_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12900_ _12900_/A _12900_/B vssd1 vssd1 vccd1 vccd1 _14141_/C sky130_fd_sc_hd__xor2_2
XFILLER_247_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13880_ _19519_/Q _13947_/A2 _13947_/B1 _13879_/X vssd1 vssd1 vccd1 vccd1 _13880_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_272_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12831_ _12936_/S _12830_/X _12746_/X vssd1 vssd1 vccd1 vccd1 _12831_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_62_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15550_ _13581_/A _15426_/B _13608_/X _15110_/X vssd1 vssd1 vccd1 vccd1 _15550_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12762_/A _12762_/B vssd1 vssd1 vccd1 vccd1 _12762_/Y sky130_fd_sc_hd__nor2_2
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _17703_/A0 _18351_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _18351_/D sky130_fd_sc_hd__mux2_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _18521_/Q _18522_/Q _18523_/Q _11711_/A vssd1 vssd1 vccd1 vccd1 _11715_/C
+ sky130_fd_sc_hd__o31a_4
XFILLER_203_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15481_/A _15481_/B vssd1 vssd1 vccd1 vccd1 _15484_/C sky130_fd_sc_hd__nand2_2
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12693_ _12613_/B _12649_/B _12729_/B vssd1 vssd1 vccd1 vccd1 _12693_/X sky130_fd_sc_hd__mux2_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _18571_/Q _17352_/A vssd1 vssd1 vccd1 vccd1 _18284_/D sky130_fd_sc_hd__and2_1
X_17220_ _19424_/Q _17256_/B vssd1 vssd1 vccd1 vccd1 _17220_/Y sky130_fd_sc_hd__nand2_1
X_11644_ _13807_/B _13761_/A _13740_/B _13810_/A vssd1 vssd1 vccd1 vccd1 _11645_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_196_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17151_ _17151_/A _17579_/A vssd1 vssd1 vccd1 vccd1 _17443_/A sky130_fd_sc_hd__nand2_1
X_14363_ _18215_/Q _17670_/A0 _14382_/S vssd1 vssd1 vccd1 vccd1 _18215_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11575_ _18267_/Q _18842_/Q _11576_/S vssd1 vssd1 vccd1 vccd1 _11575_/X sky130_fd_sc_hd__mux2_1
Xinput16 core_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_2
Xinput27 core_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
X_16102_ _16142_/A1 _16101_/Y _16149_/A vssd1 vssd1 vccd1 vccd1 _18753_/D sky130_fd_sc_hd__a21oi_1
XFILLER_156_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13314_ _12989_/Y _12994_/Y _13314_/S vssd1 vssd1 vccd1 vccd1 _13314_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput38 core_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_2
X_17082_ _17587_/A _17114_/A2 _17081_/X _17346_/A vssd1 vssd1 vccd1 vccd1 _19374_/D
+ sky130_fd_sc_hd__o211a_1
X_10526_ _10527_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _11545_/A sky130_fd_sc_hd__nor2_2
XFILLER_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput49 dout0[15] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14294_ _17712_/A0 _18153_/Q _14305_/S vssd1 vssd1 vccd1 vccd1 _18153_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16033_ _16020_/A _16056_/B _18730_/Q vssd1 vssd1 vccd1 vccd1 _16033_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13245_ _19434_/Q _12560_/B _13243_/X _13244_/X _12560_/A vssd1 vssd1 vccd1 vccd1
+ _13245_/X sky130_fd_sc_hd__o221a_1
X_10457_ _17977_/Q _11295_/A2 _11371_/B1 vssd1 vssd1 vccd1 vccd1 _10457_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13176_ _15881_/A _12506_/X _12510_/X _13175_/X vssd1 vssd1 vccd1 vccd1 _13176_/X
+ sky130_fd_sc_hd__o211a_1
X_10388_ _10386_/X _10387_/X _10785_/A vssd1 vssd1 vccd1 vccd1 _10388_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ _17836_/Q _12128_/C _17837_/Q vssd1 vssd1 vccd1 vccd1 _12129_/B sky130_fd_sc_hd__a21oi_1
XFILLER_97_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_5__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_269_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17984_ _19197_/CLK _17984_/D vssd1 vssd1 vccd1 vccd1 _17984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1840 _12428_/C1 vssd1 vssd1 vccd1 vccd1 _14179_/A sky130_fd_sc_hd__buf_2
X_16935_ _19318_/Q _17187_/B _16947_/S vssd1 vssd1 vccd1 vccd1 _16936_/B sky130_fd_sc_hd__mux2_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12058_ _12389_/A1 _12086_/A2 _12057_/X _14340_/A vssd1 vssd1 vccd1 vccd1 _17806_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_238_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1851 _16904_/A vssd1 vssd1 vccd1 vccd1 _16928_/A sky130_fd_sc_hd__clkbuf_2
Xfanout1862 fanout1863/X vssd1 vssd1 vccd1 vccd1 _15910_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1873 _16048_/A vssd1 vssd1 vccd1 vccd1 _17285_/A sky130_fd_sc_hd__buf_8
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11009_ _11481_/A _11017_/A1 _19213_/Q _11406_/B2 vssd1 vssd1 vccd1 vccd1 _11009_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout1884 fanout1905/X vssd1 vssd1 vccd1 vccd1 _12249_/A sky130_fd_sc_hd__buf_2
XFILLER_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1895 _16803_/A vssd1 vssd1 vccd1 vccd1 _16795_/A sky130_fd_sc_hd__buf_4
XFILLER_226_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16866_ _19301_/Q _17569_/A _16971_/S vssd1 vssd1 vccd1 vccd1 _16867_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18605_ _19629_/CLK _18605_/D vssd1 vssd1 vccd1 vccd1 _18605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15817_ _18609_/Q _17707_/A0 _15817_/S vssd1 vssd1 vccd1 vccd1 _18609_/D sky130_fd_sc_hd__mux2_1
XFILLER_203_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19585_ _19618_/CLK _19585_/D vssd1 vssd1 vccd1 vccd1 _19585_/Q sky130_fd_sc_hd__dfxtp_1
X_16797_ _19287_/Q _16799_/C _16796_/Y vssd1 vssd1 vccd1 vccd1 _19287_/D sky130_fd_sc_hd__a21oi_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18536_ _19592_/CLK _18536_/D vssd1 vssd1 vccd1 vccd1 _18536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _15772_/B _15748_/B vssd1 vssd1 vccd1 vccd1 _15751_/B sky130_fd_sc_hd__nor2_1
XFILLER_18_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18467_ _19646_/CLK _18467_/D vssd1 vssd1 vccd1 vccd1 _18467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15679_ _15690_/A _15677_/Y _15678_/X _15751_/A vssd1 vssd1 vccd1 vccd1 _15679_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_290 _11942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17418_ _17418_/A _17453_/B vssd1 vssd1 vccd1 vccd1 _17418_/Y sky130_fd_sc_hd__nand2_1
XFILLER_194_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18398_ _19399_/CLK _18398_/D vssd1 vssd1 vccd1 vccd1 _18398_/Q sky130_fd_sc_hd__dfxtp_4
X_17349_ _19472_/Q _17169_/B _17361_/S vssd1 vssd1 vccd1 vccd1 _17350_/B sky130_fd_sc_hd__mux2_1
XFILLER_158_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19019_ _19622_/CLK _19019_/D vssd1 vssd1 vccd1 vccd1 _19019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08984_ _08979_/Y _08983_/Y _11438_/B1 vssd1 vssd1 vccd1 vccd1 _08984_/X sky130_fd_sc_hd__a21o_1
XFILLER_244_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_164_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19546_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09605_ _09718_/S _09597_/X _09596_/X _09429_/S vssd1 vssd1 vccd1 vccd1 _09605_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_283_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09536_ _18632_/Q _18054_/Q _19073_/Q _18977_/Q _11160_/S _09857_/A1 vssd1 vssd1
+ vccd1 vccd1 _09536_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ _09463_/X _09466_/X _09690_/A vssd1 vssd1 vccd1 vccd1 _09467_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09398_ _11417_/B1 _09396_/X _09397_/X _09383_/X vssd1 vssd1 vccd1 vccd1 _09398_/X
+ sky130_fd_sc_hd__o31a_4
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ _11360_/A1 _18608_/Q _18179_/Q _11360_/B2 vssd1 vssd1 vccd1 vccd1 _11360_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10311_ _11064_/B1 _10309_/Y _10310_/X vssd1 vssd1 vccd1 vccd1 _10311_/X sky130_fd_sc_hd__o21a_1
XFILLER_285_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11291_ _11292_/A _12595_/B vssd1 vssd1 vccd1 vccd1 _11293_/A sky130_fd_sc_hd__nor2_4
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13030_ _13055_/B _13030_/B vssd1 vssd1 vccd1 vccd1 _13030_/Y sky130_fd_sc_hd__nor2_1
X_10242_ _10240_/X _10241_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _10243_/B sky130_fd_sc_hd__mux2_1
XFILLER_279_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10173_ _18265_/Q _18840_/Q _10176_/S vssd1 vssd1 vccd1 vccd1 _10173_/X sky130_fd_sc_hd__mux2_1
Xfanout1103 _15102_/Y vssd1 vssd1 vccd1 vccd1 _17559_/B sky130_fd_sc_hd__buf_4
XFILLER_121_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1114 _13874_/B vssd1 vssd1 vccd1 vccd1 _13446_/B sky130_fd_sc_hd__buf_6
Xfanout1125 _15661_/B vssd1 vssd1 vccd1 vccd1 _15793_/A2 sky130_fd_sc_hd__buf_6
XFILLER_248_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1136 _12318_/Y vssd1 vssd1 vccd1 vccd1 _15330_/A sky130_fd_sc_hd__buf_8
Xfanout1147 _09104_/X vssd1 vssd1 vccd1 vccd1 _10194_/C1 sky130_fd_sc_hd__clkbuf_16
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14981_ _18499_/Q _15011_/A2 _14980_/Y _14991_/C1 vssd1 vssd1 vccd1 vccd1 _18499_/D
+ sky130_fd_sc_hd__a211o_1
Xfanout1158 _15955_/Y vssd1 vssd1 vccd1 vccd1 _16002_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1169 _15948_/C1 vssd1 vssd1 vccd1 vccd1 _15945_/C1 sky130_fd_sc_hd__buf_4
XFILLER_75_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16720_ _19259_/Q _16723_/C _16719_/Y vssd1 vssd1 vccd1 vccd1 _19259_/D sky130_fd_sc_hd__a21oi_1
X_13932_ _13322_/Y _13916_/X _13931_/X _13915_/X _13968_/B2 vssd1 vssd1 vccd1 vccd1
+ _13932_/X sky130_fd_sc_hd__a32o_1
XFILLER_275_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16651_ _16658_/C _16651_/B vssd1 vssd1 vccd1 vccd1 _19239_/D sky130_fd_sc_hd__nor2_1
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13863_ _12704_/S _12947_/X _12953_/X _13863_/B2 vssd1 vssd1 vccd1 vccd1 _13863_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12814_ _12812_/X _12813_/X _12935_/S vssd1 vssd1 vccd1 vccd1 _12815_/A sky130_fd_sc_hd__mux2_1
X_15602_ _15638_/C _15602_/B vssd1 vssd1 vccd1 vccd1 _15602_/Y sky130_fd_sc_hd__xnor2_2
X_19370_ _19466_/CLK _19370_/D vssd1 vssd1 vccd1 vccd1 _19370_/Q sky130_fd_sc_hd__dfxtp_1
X_13794_ _13794_/A _13794_/B vssd1 vssd1 vccd1 vccd1 _14151_/B sky130_fd_sc_hd__xnor2_4
X_16582_ _16615_/A0 _19186_/Q _16585_/S vssd1 vssd1 vccd1 vccd1 _19186_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18321_ _19600_/CLK _18321_/D vssd1 vssd1 vccd1 vccd1 _18321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15533_ _18581_/Q _15561_/C vssd1 vssd1 vccd1 vccd1 _15581_/C sky130_fd_sc_hd__and2_1
X_12745_ _13314_/S _12746_/B vssd1 vssd1 vccd1 vccd1 _12745_/X sky130_fd_sc_hd__or2_4
XFILLER_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _19147_/CLK _18252_/D vssd1 vssd1 vccd1 vccd1 _18252_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ _15464_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _15464_/X sky130_fd_sc_hd__or2_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _11136_/Y _12596_/B _12733_/S vssd1 vssd1 vccd1 vccd1 _12676_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14415_ _16622_/A0 _18266_/Q _14415_/S vssd1 vssd1 vccd1 vccd1 _18266_/D sky130_fd_sc_hd__mux2_1
X_17203_ _19419_/Q fanout533/X _17202_/Y _17119_/B vssd1 vssd1 vccd1 vccd1 _17204_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_11627_ _11628_/A _13962_/A vssd1 vssd1 vccd1 vccd1 _11627_/Y sky130_fd_sc_hd__nor2_4
X_18183_ _19631_/CLK _18183_/D vssd1 vssd1 vccd1 vccd1 _18183_/Q sky130_fd_sc_hd__dfxtp_1
X_15395_ _15376_/A _15376_/B _15373_/A vssd1 vssd1 vccd1 vccd1 _15399_/A sky130_fd_sc_hd__o21ai_4
XFILLER_128_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14346_ _14487_/A _14346_/B vssd1 vssd1 vccd1 vccd1 _18201_/D sky130_fd_sc_hd__nor2_1
X_17134_ _19396_/Q fanout534/X _17413_/A _17212_/B2 vssd1 vssd1 vccd1 vccd1 _17135_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_184_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11558_ _17983_/Q _16820_/A3 _08947_/X _17951_/Q _11557_/Y vssd1 vssd1 vccd1 vccd1
+ _11558_/X sky130_fd_sc_hd__a221o_4
XFILLER_183_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17065_ _19366_/Q _17077_/B vssd1 vssd1 vccd1 vccd1 _17065_/X sky130_fd_sc_hd__or2_1
XFILLER_156_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ _10662_/A1 _19220_/Q _19188_/Q _10656_/S _08899_/A vssd1 vssd1 vccd1 vccd1
+ _10509_/X sky130_fd_sc_hd__a221o_1
XFILLER_144_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14277_ _17695_/A0 _18136_/Q _14277_/S vssd1 vssd1 vccd1 vccd1 _18136_/D sky130_fd_sc_hd__mux2_1
XFILLER_195_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11489_ _17900_/Q _11490_/B _11489_/B1 _11488_/Y vssd1 vssd1 vccd1 vccd1 _12625_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_143_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16016_ _18723_/Q _16016_/A2 _16147_/A2 _18772_/Q _16018_/C1 vssd1 vssd1 vccd1 vccd1
+ _16016_/X sky130_fd_sc_hd__a221o_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ _12875_/X _12888_/Y _13354_/A vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _18109_/Q _18108_/Q _13159_/C vssd1 vssd1 vccd1 vccd1 _13201_/B sky130_fd_sc_hd__and3_1
XFILLER_285_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _17975_/CLK _17967_/D vssd1 vssd1 vccd1 vccd1 _17967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1670 _09958_/C1 vssd1 vssd1 vccd1 vccd1 _08895_/A sky130_fd_sc_hd__buf_12
X_16918_ _16970_/A1 _17938_/Q _16917_/X vssd1 vssd1 vccd1 vccd1 _17175_/B sky130_fd_sc_hd__o21a_4
XFILLER_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1681 _09854_/A vssd1 vssd1 vccd1 vccd1 _11566_/A1 sky130_fd_sc_hd__buf_4
Xfanout1692 _11404_/A1 vssd1 vssd1 vccd1 vccd1 _11469_/A1 sky130_fd_sc_hd__buf_6
X_17898_ _18201_/CLK _17898_/D vssd1 vssd1 vccd1 vccd1 _17898_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_265_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_19637_ _19637_/CLK _19637_/D vssd1 vssd1 vccd1 vccd1 _19637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16849_ _16850_/B vssd1 vssd1 vccd1 vccd1 _17123_/B sky130_fd_sc_hd__clkinv_4
XFILLER_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19568_ _19600_/CLK _19568_/D vssd1 vssd1 vccd1 vccd1 _19568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09321_ _09908_/A1 _09232_/A _09320_/X _09908_/B1 _18397_/Q vssd1 vssd1 vccd1 vccd1
+ _09986_/C sky130_fd_sc_hd__o32a_2
X_18519_ _19291_/CLK _18519_/D vssd1 vssd1 vccd1 vccd1 _18519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19499_ _19531_/CLK _19499_/D vssd1 vssd1 vccd1 vccd1 _19499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _18541_/Q _18416_/Q _09252_/S vssd1 vssd1 vccd1 vccd1 _09252_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09183_ _11389_/A1 _18214_/Q _09181_/S _18949_/Q _11001_/C1 vssd1 vssd1 vccd1 vccd1
+ _09183_/X sky130_fd_sc_hd__o221a_1
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput206 localMemory_wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput217 localMemory_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input217/X sky130_fd_sc_hd__buf_8
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput228 localMemory_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 input228/X sky130_fd_sc_hd__clkbuf_16
X_08967_ _08965_/X _08966_/X _08967_/S vssd1 vssd1 vccd1 vccd1 _08967_/X sky130_fd_sc_hd__mux2_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput239 localMemory_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 input239/X sky130_fd_sc_hd__buf_12
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08898_ _17906_/Q _09062_/B vssd1 vssd1 vccd1 vccd1 _08898_/Y sky130_fd_sc_hd__nand2_8
XFILLER_257_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _18831_/Q _11300_/B vssd1 vssd1 vccd1 vccd1 _10860_/X sky130_fd_sc_hd__or2_1
XFILLER_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09519_ _09976_/A1 _09517_/X _09518_/X _11198_/S vssd1 vssd1 vccd1 vccd1 _09519_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10791_ _11332_/B1 _10790_/X _11800_/B vssd1 vssd1 vccd1 vccd1 _10791_/X sky130_fd_sc_hd__o21a_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _19328_/Q _12524_/Y _12529_/Y _19456_/Q _12516_/Y vssd1 vssd1 vccd1 vccd1
+ _12530_/X sky130_fd_sc_hd__a221o_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19126_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ _12461_/A _13462_/A vssd1 vssd1 vccd1 vccd1 _12461_/Y sky130_fd_sc_hd__nand2_4
XFILLER_185_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14200_ _18711_/Q _18098_/Q _14200_/S vssd1 vssd1 vccd1 vccd1 _14201_/B sky130_fd_sc_hd__mux2_1
XFILLER_138_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11412_ _17901_/Q _11490_/B _11489_/B1 _11411_/Y vssd1 vssd1 vccd1 vccd1 _12597_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_137_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15180_ _15200_/B _15179_/X _15113_/Y vssd1 vssd1 vccd1 vccd1 _15192_/B sky130_fd_sc_hd__o21a_1
X_12392_ _08896_/A _12430_/A _12391_/Y _14001_/C1 vssd1 vssd1 vccd1 vccd1 _17905_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_193_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14131_ _16548_/A0 _18070_/Q _14131_/S vssd1 vssd1 vccd1 vccd1 _18070_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11343_ _11358_/A _11338_/X _11342_/X vssd1 vssd1 vccd1 vccd1 _11343_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_192_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ _16314_/A0 _18004_/Q _14073_/S vssd1 vssd1 vccd1 vccd1 _18004_/D sky130_fd_sc_hd__mux2_1
X_11274_ _18641_/Q _18063_/Q _19082_/Q _18986_/Q _11617_/S _11274_/S1 vssd1 vssd1
+ vccd1 vccd1 _11275_/B sky130_fd_sc_hd__mux4_1
XFILLER_153_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13013_ _19301_/Q _13952_/A2 _12551_/Y vssd1 vssd1 vccd1 vccd1 _13013_/X sky130_fd_sc_hd__a21o_1
X_10225_ _10223_/X _10224_/X _10225_/S vssd1 vssd1 vccd1 vccd1 _10225_/X sky130_fd_sc_hd__mux2_1
X_18870_ _18902_/CLK _18870_/D vssd1 vssd1 vccd1 vccd1 _18870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17821_ _19490_/CLK _17821_/D vssd1 vssd1 vccd1 vccd1 _17821_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10156_ _13917_/A vssd1 vssd1 vccd1 vccd1 _10156_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17752_ _18652_/Q vssd1 vssd1 vccd1 vccd1 _18652_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_248_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10087_ _11143_/A1 _10086_/Y _10082_/X vssd1 vssd1 vccd1 vccd1 _10087_/X sky130_fd_sc_hd__o21a_1
X_14964_ _14962_/X _14963_/X _14964_/B1 vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__a21o_1
XFILLER_75_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16703_ _19253_/Q _16708_/D _19254_/Q vssd1 vssd1 vccd1 vccd1 _16705_/B sky130_fd_sc_hd__a21oi_1
XFILLER_263_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13915_ _13966_/C1 _13911_/Y _13914_/X _13910_/X vssd1 vssd1 vccd1 vccd1 _13915_/X
+ sky130_fd_sc_hd__a31o_1
X_17683_ _17683_/A0 _19610_/Q _17690_/S vssd1 vssd1 vccd1 vccd1 _19610_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14895_ _15835_/B _16078_/C _11715_/B vssd1 vssd1 vccd1 vccd1 _14895_/X sky130_fd_sc_hd__a21bo_1
XFILLER_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19422_ _19552_/CLK _19422_/D vssd1 vssd1 vccd1 vccd1 _19422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16634_ _16752_/A _16634_/B _16677_/A vssd1 vssd1 vccd1 vccd1 _19233_/D sky130_fd_sc_hd__nor3_1
X_13846_ _17851_/Q _13846_/B vssd1 vssd1 vccd1 vccd1 _13846_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19353_ _19481_/CLK _19353_/D vssd1 vssd1 vccd1 vccd1 _19353_/Q sky130_fd_sc_hd__dfxtp_1
X_13777_ _19258_/Q _13943_/A2 _13943_/B1 _19290_/Q vssd1 vssd1 vccd1 vccd1 _13777_/X
+ sky130_fd_sc_hd__a22o_1
X_16565_ _17665_/A0 _19169_/Q _16586_/S vssd1 vssd1 vccd1 vccd1 _19169_/D sky130_fd_sc_hd__mux2_1
XFILLER_222_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10989_ _17938_/Q _11451_/A2 _10988_/Y _11451_/B2 vssd1 vssd1 vccd1 vccd1 _10989_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18304_ _19453_/CLK _18304_/D vssd1 vssd1 vccd1 vccd1 _18304_/Q sky130_fd_sc_hd__dfxtp_1
X_15516_ _15537_/B1 _15514_/Y _15515_/Y _15751_/A vssd1 vssd1 vccd1 vccd1 _15516_/X
+ sky130_fd_sc_hd__a211o_1
X_19284_ _19295_/CLK _19284_/D vssd1 vssd1 vccd1 vccd1 _19284_/Q sky130_fd_sc_hd__dfxtp_1
X_12728_ _12600_/B _12639_/B _12733_/S vssd1 vssd1 vccd1 vccd1 _12728_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16496_ _16529_/A0 _19102_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _19102_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18235_ _19134_/CLK _18235_/D vssd1 vssd1 vccd1 vccd1 _18235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12659_ _11633_/Y _12658_/Y _12657_/Y vssd1 vssd1 vccd1 vccd1 _12659_/Y sky130_fd_sc_hd__o21ai_2
X_15447_ _18577_/Q _15447_/B vssd1 vssd1 vccd1 vccd1 _15447_/Y sky130_fd_sc_hd__nor2_1
XFILLER_276_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18166_ _19619_/CLK _18166_/D vssd1 vssd1 vccd1 vccd1 _18166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15378_ _17389_/B1 _15377_/X _15499_/B1 vssd1 vssd1 vccd1 vccd1 _15378_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17117_ _17157_/A _17117_/B vssd1 vssd1 vccd1 vccd1 _17394_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ _18186_/Q _17713_/A0 _14339_/S vssd1 vssd1 vccd1 vccd1 _18186_/D sky130_fd_sc_hd__mux2_1
X_18097_ _18713_/CLK _18097_/D vssd1 vssd1 vccd1 vccd1 _18097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17048_ _17048_/A _17555_/B vssd1 vssd1 vccd1 vccd1 _17591_/D sky130_fd_sc_hd__or2_4
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout907 _16426_/X vssd1 vssd1 vccd1 vccd1 _16458_/S sky130_fd_sc_hd__buf_8
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _10742_/A1 _09868_/X _09869_/X _11607_/S vssd1 vssd1 vccd1 vccd1 _09870_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout918 _16278_/S vssd1 vssd1 vccd1 vccd1 _16288_/S sky130_fd_sc_hd__buf_12
XFILLER_258_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 _17475_/B1 vssd1 vssd1 vccd1 vccd1 _17543_/B1 sky130_fd_sc_hd__buf_2
XFILLER_97_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08821_ _19295_/Q vssd1 vssd1 vccd1 vccd1 _08821_/Y sky130_fd_sc_hd__inv_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18999_ _19138_/CLK _18999_/D vssd1 vssd1 vccd1 vccd1 _18999_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09304_ _19108_/Q _19140_/Q _09306_/S vssd1 vssd1 vccd1 vccd1 _09304_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09235_ input115/X input150/X _09657_/S vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__mux2_4
XFILLER_210_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09166_ _10169_/S _09164_/X _09165_/X vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__a21o_1
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09097_ _14074_/B _09683_/A vssd1 vssd1 vccd1 vccd1 _09097_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_134_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10010_ _18594_/Q _18165_/Q _10840_/S vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__mux2_1
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ _11566_/A1 _18204_/Q _11226_/S _18939_/Q _11569_/S1 vssd1 vssd1 vccd1 vccd1
+ _09999_/X sky130_fd_sc_hd__o221a_1
XFILLER_131_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ _18507_/Q _11720_/X _11911_/X _11968_/B2 vssd1 vssd1 vccd1 vccd1 _11961_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10912_ _10912_/A _10912_/B vssd1 vssd1 vccd1 vccd1 _10912_/Y sky130_fd_sc_hd__nor2_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _11541_/B _13962_/B _13153_/X _12732_/S _13699_/Y vssd1 vssd1 vccd1 vccd1
+ _13700_/X sky130_fd_sc_hd__o221a_1
XFILLER_245_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _14688_/B _14680_/B _14680_/C _14672_/C vssd1 vssd1 vccd1 vccd1 _14993_/S
+ sky130_fd_sc_hd__or4b_4
XFILLER_205_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11892_ _11819_/X _11875_/A _11901_/B _11854_/X vssd1 vssd1 vccd1 vccd1 _11892_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13631_ _19445_/Q _13655_/A2 _13629_/X _13630_/X _13655_/C1 vssd1 vssd1 vccd1 vccd1
+ _13631_/X sky130_fd_sc_hd__o221a_1
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10843_ _11584_/A1 _19151_/Q _11581_/S _19119_/Q _11562_/S vssd1 vssd1 vccd1 vccd1
+ _10843_/X sky130_fd_sc_hd__o221a_1
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16350_ _18962_/Q _17682_/A0 _16358_/S vssd1 vssd1 vccd1 vccd1 _18962_/D sky130_fd_sc_hd__mux2_1
X_13562_ _13757_/A _14012_/B _13548_/X vssd1 vssd1 vccd1 vccd1 _13562_/Y sky130_fd_sc_hd__o21ai_1
X_10774_ _11584_/C1 _10771_/X _10773_/X vssd1 vssd1 vccd1 vccd1 _10774_/X sky130_fd_sc_hd__a21o_1
XFILLER_185_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12513_ _12499_/A _12513_/B vssd1 vssd1 vccd1 vccd1 _12514_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15301_ _17129_/A _15300_/X _15424_/C1 vssd1 vssd1 vccd1 vccd1 _15301_/X sky130_fd_sc_hd__a21o_1
XFILLER_200_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16281_ _17712_/A0 _18895_/Q _16292_/S vssd1 vssd1 vccd1 vccd1 _18895_/D sky130_fd_sc_hd__mux2_1
X_13493_ _17840_/Q _13744_/A2 _13744_/B1 _17872_/Q vssd1 vssd1 vccd1 vccd1 _13493_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18020_ _19622_/CLK _18020_/D vssd1 vssd1 vccd1 vccd1 _18020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12444_ _12445_/A _12445_/B vssd1 vssd1 vccd1 vccd1 _12444_/X sky130_fd_sc_hd__and2_4
X_15232_ _19461_/Q _19395_/Q _15231_/X vssd1 vssd1 vccd1 vccd1 _15233_/B sky130_fd_sc_hd__o21ai_4
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15163_ _15163_/A _15163_/B vssd1 vssd1 vccd1 vccd1 _15163_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12375_ _18385_/Q _12429_/B1 _09653_/B _08858_/A vssd1 vssd1 vccd1 vccd1 _12376_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_5_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14114_ _16465_/A0 _18053_/Q _14131_/S vssd1 vssd1 vccd1 vccd1 _18053_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11326_ _11572_/A1 _18147_/Q _18793_/Q _11325_/S vssd1 vssd1 vccd1 vccd1 _11326_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15094_ _19376_/Q _15086_/B input171/X _15086_/X vssd1 vssd1 vccd1 vccd1 _15094_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_153_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14045_ _16595_/A0 _17987_/Q _14073_/S vssd1 vssd1 vccd1 vccd1 _17987_/D sky130_fd_sc_hd__mux2_1
X_18922_ _19640_/CLK _18922_/D vssd1 vssd1 vccd1 vccd1 _18922_/Q sky130_fd_sc_hd__dfxtp_1
X_11257_ _09859_/A _17641_/A0 _11256_/X _11257_/C1 vssd1 vssd1 vccd1 vccd1 _11832_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_140_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10208_ _10200_/S _10206_/X _10207_/X _10356_/C1 vssd1 vssd1 vccd1 vccd1 _10208_/X
+ sky130_fd_sc_hd__a211o_1
X_18853_ _19203_/CLK _18853_/D vssd1 vssd1 vccd1 vccd1 _18853_/Q sky130_fd_sc_hd__dfxtp_1
X_11188_ _18642_/Q _18064_/Q _19083_/Q _18987_/Q _09885_/S _11274_/S1 vssd1 vssd1
+ vccd1 vccd1 _11189_/B sky130_fd_sc_hd__mux4_1
XFILLER_67_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17804_ _19650_/CLK _17804_/D vssd1 vssd1 vccd1 vccd1 _17804_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10139_ _10219_/A1 _19225_/Q _19193_/Q _10215_/S _10293_/B1 vssd1 vssd1 vccd1 vccd1
+ _10139_/X sky130_fd_sc_hd__a221o_1
X_18784_ _18902_/CLK _18784_/D vssd1 vssd1 vccd1 vccd1 _18784_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _18713_/Q _16002_/A2 _16004_/B1 _18762_/Q _16004_/C1 vssd1 vssd1 vccd1 vccd1
+ _15996_/X sky130_fd_sc_hd__a221o_1
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17735_ _18635_/Q vssd1 vssd1 vccd1 vccd1 _18635_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14947_ input60/X input95/X _14947_/S vssd1 vssd1 vccd1 vccd1 _14948_/A sky130_fd_sc_hd__mux2_2
XFILLER_209_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17666_ _17666_/A0 _19593_/Q _17687_/S vssd1 vssd1 vccd1 vccd1 _19593_/D sky130_fd_sc_hd__mux2_1
X_14878_ _14696_/A _18271_/Q _14877_/Y _14918_/B1 vssd1 vssd1 vccd1 vccd1 _14878_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_78_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19405_ _19530_/CLK _19405_/D vssd1 vssd1 vccd1 vccd1 _19405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16617_ _16617_/A0 _19220_/Q _16618_/S vssd1 vssd1 vccd1 vccd1 _19220_/D sky130_fd_sc_hd__mux2_1
XFILLER_211_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13829_ _19323_/Q _13952_/A2 _13854_/B1 _13822_/X _13828_/X vssd1 vssd1 vccd1 vccd1
+ _13829_/Y sky130_fd_sc_hd__a2111oi_2
XFILLER_211_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17597_ _19378_/Q _15086_/B input179/X _17592_/X _17623_/B1 vssd1 vssd1 vccd1 vccd1
+ _17597_/X sky130_fd_sc_hd__a41o_1
X_19336_ _19464_/CLK _19336_/D vssd1 vssd1 vccd1 vccd1 _19336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16548_ _16548_/A0 _19153_/Q _16548_/S vssd1 vssd1 vccd1 vccd1 _19153_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19267_ _19268_/CLK _19267_/D vssd1 vssd1 vccd1 vccd1 _19267_/Q sky130_fd_sc_hd__dfxtp_1
X_16479_ _17711_/A0 _19086_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _19086_/D sky130_fd_sc_hd__mux2_1
X_09020_ _09043_/A _09031_/S vssd1 vssd1 vccd1 vccd1 _09039_/B sky130_fd_sc_hd__nand2_4
X_18218_ _19600_/CLK _18218_/D vssd1 vssd1 vccd1 vccd1 _18218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19198_ _19621_/CLK _19198_/D vssd1 vssd1 vccd1 vccd1 _19198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18149_ _19211_/CLK _18149_/D vssd1 vssd1 vccd1 vccd1 _18149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09922_ _09683_/A _09920_/X _09921_/X _10996_/B1 _09919_/X vssd1 vssd1 vccd1 vccd1
+ _09922_/X sky130_fd_sc_hd__o311a_1
Xfanout704 _12544_/Y vssd1 vssd1 vccd1 vccd1 _13425_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout715 _12919_/A2 vssd1 vssd1 vccd1 vccd1 _13945_/A2 sky130_fd_sc_hd__buf_4
Xfanout726 _12495_/Y vssd1 vssd1 vccd1 vccd1 _13942_/A2 sky130_fd_sc_hd__buf_6
Xfanout737 _16507_/A0 vssd1 vssd1 vccd1 vccd1 _17706_/A0 sky130_fd_sc_hd__clkbuf_4
X_09853_ _09850_/X _09852_/X _09853_/S vssd1 vssd1 vccd1 vccd1 _09853_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout748 _09779_/X vssd1 vssd1 vccd1 vccd1 _13263_/A sky130_fd_sc_hd__buf_6
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout759 _16470_/A0 vssd1 vssd1 vccd1 vccd1 _17669_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09784_ _18239_/Q _18814_/Q _09797_/S vssd1 vssd1 vccd1 vccd1 _09784_/X sky130_fd_sc_hd__mux2_1
XFILLER_258_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_108 _11732_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_119 _11820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09218_ _19077_/Q _18981_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _09218_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10490_ _17913_/Q _11135_/S _11181_/B1 _10489_/Y vssd1 vssd1 vccd1 vccd1 _10527_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09149_ input116/X input152/X _09657_/S vssd1 vssd1 vccd1 vccd1 _09149_/X sky130_fd_sc_hd__mux2_8
XFILLER_182_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _17848_/Q _17849_/Q _12160_/C vssd1 vssd1 vccd1 vccd1 _12162_/B sky130_fd_sc_hd__and3_1
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11111_ _18643_/Q _18065_/Q _19084_/Q _18988_/Q _11609_/S _11622_/A1 vssd1 vssd1
+ vccd1 vccd1 _11112_/B sky130_fd_sc_hd__mux4_1
X_12091_ _12107_/A _17823_/Q vssd1 vssd1 vccd1 vccd1 _17823_/D sky130_fd_sc_hd__nor2_1
XFILLER_146_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _11040_/X _11041_/X _11507_/S vssd1 vssd1 vccd1 vccd1 _11042_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _15853_/A _15955_/B vssd1 vssd1 vccd1 vccd1 _15850_/X sky130_fd_sc_hd__and2_1
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _18112_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14801_/X sky130_fd_sc_hd__or2_1
XFILLER_18_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _19486_/Q _15780_/Y _15781_/S vssd1 vssd1 vccd1 vccd1 _15781_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _12684_/Y _12727_/X _13089_/A vssd1 vssd1 vccd1 vccd1 _12994_/A sky130_fd_sc_hd__mux2_2
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _13807_/B _17520_/A2 _17543_/B1 _17816_/Q _17550_/A vssd1 vssd1 vccd1 vccd1
+ _17520_/X sky130_fd_sc_hd__a221o_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _17794_/Q _14982_/B vssd1 vssd1 vccd1 vccd1 _14732_/X sky130_fd_sc_hd__or2_1
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ _11944_/A1 _11878_/B _11878_/C _11959_/A2 input231/X vssd1 vssd1 vccd1 vccd1
+ _11944_/X sky130_fd_sc_hd__a32o_4
XFILLER_245_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17451_ _18574_/Q _17527_/A1 _17546_/A2 vssd1 vssd1 vccd1 vccd1 _17451_/X sky130_fd_sc_hd__o21a_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14663_ _17722_/A0 _18469_/Q _14663_/S vssd1 vssd1 vccd1 vccd1 _18469_/D sky130_fd_sc_hd__mux2_1
X_11875_ _11875_/A _11901_/B vssd1 vssd1 vccd1 vccd1 _11875_/Y sky130_fd_sc_hd__nand2_8
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _17667_/A0 _19011_/Q _16424_/S vssd1 vssd1 vccd1 vccd1 _19011_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10826_ _10819_/X _10825_/X _10809_/X vssd1 vssd1 vccd1 vccd1 _10826_/Y sky130_fd_sc_hd__o21ai_4
X_13614_ _13622_/B _13961_/A vssd1 vssd1 vccd1 vccd1 _13614_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17382_ _17382_/A _17382_/B vssd1 vssd1 vccd1 vccd1 _17386_/B sky130_fd_sc_hd__nor2_1
X_14594_ _14522_/Y _08884_/X input9/X _14525_/A vssd1 vssd1 vccd1 vccd1 _14594_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19121_ _19602_/CLK _19121_/D vssd1 vssd1 vccd1 vccd1 _19121_/Q sky130_fd_sc_hd__dfxtp_1
X_16333_ _18945_/Q _16532_/A0 _16352_/S vssd1 vssd1 vccd1 vccd1 _18945_/D sky130_fd_sc_hd__mux2_1
X_10757_ _11556_/C _10757_/B vssd1 vssd1 vccd1 vccd1 _10757_/Y sky130_fd_sc_hd__nor2_1
X_13545_ _13545_/A _13545_/B vssd1 vssd1 vccd1 vccd1 _13545_/X sky130_fd_sc_hd__or2_1
XFILLER_41_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19052_ _19621_/CLK _19052_/D vssd1 vssd1 vccd1 vccd1 _19052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13476_ _13937_/A _13476_/B vssd1 vssd1 vccd1 vccd1 _13476_/X sky130_fd_sc_hd__or2_1
X_16264_ _17662_/A0 _18878_/Q _16278_/S vssd1 vssd1 vccd1 vccd1 _18878_/D sky130_fd_sc_hd__mux2_1
X_10688_ _11173_/S _10687_/X _10686_/X vssd1 vssd1 vccd1 vccd1 _10688_/X sky130_fd_sc_hd__o21a_1
X_18003_ _19573_/CLK _18003_/D vssd1 vssd1 vccd1 vccd1 _18003_/Q sky130_fd_sc_hd__dfxtp_1
X_12427_ _12427_/A _12427_/B vssd1 vssd1 vccd1 vccd1 _12427_/Y sky130_fd_sc_hd__nand2_1
X_15215_ _15304_/A1 _13056_/X _15285_/A3 _15214_/X vssd1 vssd1 vccd1 vccd1 _15215_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16195_ _17692_/A0 _18811_/Q _16212_/S vssd1 vssd1 vccd1 vccd1 _18811_/D sky130_fd_sc_hd__mux2_1
Xoutput307 _11755_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[11] sky130_fd_sc_hd__buf_4
XFILLER_236_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12358_ _12421_/A _12358_/B vssd1 vssd1 vccd1 vccd1 _12358_/Y sky130_fd_sc_hd__nand2_1
Xoutput318 _11765_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[21] sky130_fd_sc_hd__buf_4
X_15146_ _17382_/A _15139_/X _15140_/Y _15145_/X _15351_/A2 vssd1 vssd1 vccd1 vccd1
+ _15147_/B sky130_fd_sc_hd__o311a_1
XFILLER_141_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput329 _11744_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[6] sky130_fd_sc_hd__buf_4
XFILLER_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11309_ _18030_/Q _17998_/Q _11309_/S vssd1 vssd1 vccd1 vccd1 _11309_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15077_ _18561_/Q _17688_/A0 _15078_/S vssd1 vssd1 vccd1 vccd1 _18561_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12289_ _18087_/Q _12277_/B _14934_/C _18510_/Q vssd1 vssd1 vccd1 vccd1 _14682_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_142_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18905_ _19193_/CLK _18905_/D vssd1 vssd1 vccd1 vccd1 _18905_/Q sky130_fd_sc_hd__dfxtp_1
X_14028_ _14028_/A _14028_/B vssd1 vssd1 vccd1 vccd1 _14028_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18836_ _19643_/CLK _18836_/D vssd1 vssd1 vccd1 vccd1 _18836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18767_ _18772_/CLK _18767_/D vssd1 vssd1 vccd1 vccd1 _18767_/Q sky130_fd_sc_hd__dfxtp_1
X_15979_ _18705_/Q _16019_/A2 _15978_/X _16972_/A vssd1 vssd1 vccd1 vccd1 _18705_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17718_ _17718_/A0 _19644_/Q _17718_/S vssd1 vssd1 vccd1 vccd1 _19644_/D sky130_fd_sc_hd__mux2_1
X_18698_ _19304_/CLK _18698_/D vssd1 vssd1 vccd1 vccd1 _18698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17649_ _17682_/A0 _19577_/Q _17657_/S vssd1 vssd1 vccd1 vccd1 _19577_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_189_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19154_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19319_ _19319_/CLK _19319_/D vssd1 vssd1 vccd1 vccd1 _19319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_118_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19295_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09003_ _11691_/B1 _09652_/A _09002_/X _11692_/A1 _18388_/Q vssd1 vssd1 vccd1 vccd1
+ _11217_/C sky130_fd_sc_hd__o32a_1
XFILLER_164_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout501 _11959_/B2 vssd1 vssd1 vccd1 vccd1 _11939_/A1 sky130_fd_sc_hd__buf_6
XFILLER_259_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09905_ _09903_/B _09903_/C _09903_/D _09028_/B vssd1 vssd1 vccd1 vccd1 _09905_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout512 _17499_/A2 vssd1 vssd1 vccd1 vccd1 _17462_/B sky130_fd_sc_hd__clkbuf_8
Xfanout523 _15447_/B vssd1 vssd1 vccd1 vccd1 _15351_/A2 sky130_fd_sc_hd__buf_6
XFILLER_116_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout534 fanout536/X vssd1 vssd1 vccd1 vccd1 fanout534/X sky130_fd_sc_hd__buf_6
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout545 _15476_/A1 vssd1 vssd1 vccd1 vccd1 _17129_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_247_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout556 _15122_/Y vssd1 vssd1 vccd1 vccd1 _17151_/A sky130_fd_sc_hd__clkbuf_4
Xfanout567 _15124_/X vssd1 vssd1 vccd1 vccd1 _15731_/B1 sky130_fd_sc_hd__buf_8
X_09836_ _11157_/A1 _19197_/Q _19165_/Q _11147_/S vssd1 vssd1 vccd1 vccd1 _09836_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout578 _12338_/Y vssd1 vssd1 vccd1 vccd1 _12379_/A sky130_fd_sc_hd__buf_2
XFILLER_112_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout589 _12073_/B vssd1 vssd1 vccd1 vccd1 _12085_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_47_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09767_ _09764_/X _09766_/X _10399_/A vssd1 vssd1 vccd1 vccd1 _09768_/B sky130_fd_sc_hd__a21oi_1
XFILLER_215_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09698_ _09696_/X _09697_/Y _09946_/B1 vssd1 vssd1 vccd1 vccd1 _09735_/A sky130_fd_sc_hd__a21oi_4
XFILLER_215_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _11845_/B _11887_/B1 _11659_/X _11846_/A vssd1 vssd1 vccd1 vccd1 _15120_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_186_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _18462_/Q _18363_/Q _10619_/S vssd1 vssd1 vccd1 vccd1 _10611_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11591_ _10532_/A _17723_/A0 _11590_/Y _11800_/B vssd1 vssd1 vccd1 vccd1 _11591_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_167_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13330_ _13938_/A _13330_/B vssd1 vssd1 vccd1 vccd1 _13330_/Y sky130_fd_sc_hd__nand2_1
X_10542_ _18618_/Q _18189_/Q _10619_/S vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13261_ _13261_/A _13261_/B vssd1 vssd1 vccd1 vccd1 _13261_/X sky130_fd_sc_hd__xor2_1
X_10473_ _10623_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10473_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ _17868_/Q _12210_/B _12211_/Y vssd1 vssd1 vccd1 vccd1 _17868_/D sky130_fd_sc_hd__o21a_1
X_15000_ _14996_/Y _14999_/X _15010_/B1 vssd1 vssd1 vccd1 vccd1 _15000_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13192_ _12807_/X _12827_/X _13354_/A vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12143_ _17842_/Q _12144_/C _17843_/Q vssd1 vssd1 vccd1 vccd1 _12145_/B sky130_fd_sc_hd__a21oi_1
XFILLER_269_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_4__f_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_4__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16951_ _19322_/Q _17199_/B _16971_/S vssd1 vssd1 vccd1 vccd1 _16952_/B sky130_fd_sc_hd__mux2_1
X_12074_ _11252_/S _12086_/A2 _12073_/X _14340_/A vssd1 vssd1 vccd1 vccd1 _17814_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_278_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15902_ _15902_/A _15905_/B _15905_/C vssd1 vssd1 vccd1 vccd1 _15902_/X sky130_fd_sc_hd__and3_1
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11025_ _11103_/A _11845_/A vssd1 vssd1 vccd1 vccd1 _11025_/Y sky130_fd_sc_hd__nor2_1
X_16882_ _16898_/A1 _17929_/Q _16881_/X vssd1 vssd1 vccd1 vccd1 _17577_/A sky130_fd_sc_hd__o21a_4
XFILLER_103_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18621_ _19608_/CLK _18621_/D vssd1 vssd1 vccd1 vccd1 _18621_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _18625_/Q _16292_/A0 _15833_/S vssd1 vssd1 vccd1 vccd1 _18625_/D sky130_fd_sc_hd__mux2_1
XFILLER_237_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _19575_/CLK _18552_/D vssd1 vssd1 vccd1 vccd1 _18552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _15764_/A _15765_/B vssd1 vssd1 vccd1 vccd1 _15766_/A sky130_fd_sc_hd__nand2_1
X_12976_ _17859_/Q _13945_/A2 _12965_/X _13303_/B2 _13952_/B1 vssd1 vssd1 vccd1 vccd1
+ _12977_/B sky130_fd_sc_hd__a221o_1
XFILLER_205_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _17503_/A _17523_/B vssd1 vssd1 vccd1 vccd1 _17503_/Y sky130_fd_sc_hd__nand2_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _14964_/B1 _14713_/X _14714_/Y _14690_/Y vssd1 vssd1 vccd1 vccd1 _14715_/X
+ sky130_fd_sc_hd__o211a_1
X_18483_ _19323_/CLK _18483_/D vssd1 vssd1 vccd1 vccd1 _18483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _11959_/B2 _11802_/B _11935_/B1 input244/X vssd1 vssd1 vccd1 vccd1 _11927_/X
+ sky130_fd_sc_hd__a22o_4
X_15695_ _15693_/Y _15695_/B vssd1 vssd1 vccd1 vccd1 _15696_/B sky130_fd_sc_hd__and2b_1
XFILLER_45_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_450 _14026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_461 _18373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_472 input205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17434_ _19498_/Q _17462_/B _17432_/X _17433_/Y _17338_/A vssd1 vssd1 vccd1 vccd1
+ _19498_/D sky130_fd_sc_hd__o221a_1
X_14646_ _17705_/A0 _18452_/Q _14663_/S vssd1 vssd1 vccd1 vccd1 _18452_/D sky130_fd_sc_hd__mux2_1
XANTENNA_483 input242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_494 _18106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11858_ _11859_/A _11858_/B vssd1 vssd1 vccd1 vccd1 _11863_/B sky130_fd_sc_hd__or2_1
XFILLER_159_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_19 _14929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10809_ _11131_/A _10803_/X _10806_/X _10808_/X _11623_/A1 vssd1 vssd1 vccd1 vccd1
+ _10809_/X sky130_fd_sc_hd__a311o_4
X_17365_ _19480_/Q _17193_/B _17379_/S vssd1 vssd1 vccd1 vccd1 _17366_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11789_ _11799_/A _11799_/B _11846_/B vssd1 vssd1 vccd1 vccd1 _11789_/X sky130_fd_sc_hd__and3_1
X_14577_ _18397_/Q _14589_/A2 _14589_/B1 input26/X vssd1 vssd1 vccd1 vccd1 _14578_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19104_ _19608_/CLK _19104_/D vssd1 vssd1 vccd1 vccd1 _19104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16316_ _17714_/A0 _18929_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _18929_/D sky130_fd_sc_hd__mux2_1
X_13528_ _13929_/A1 _13527_/X _13515_/Y vssd1 vssd1 vccd1 vccd1 _13528_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17296_ _18126_/Q _15717_/B2 _17517_/A _17289_/B vssd1 vssd1 vccd1 vccd1 _17296_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_146_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19035_ _19618_/CLK _19035_/D vssd1 vssd1 vccd1 vccd1 _19035_/Q sky130_fd_sc_hd__dfxtp_1
X_16247_ _16611_/A0 _18862_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _18862_/D sky130_fd_sc_hd__mux2_1
X_13459_ _14006_/B vssd1 vssd1 vccd1 vccd1 _13459_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16178_ _16608_/A0 _18795_/Q _16189_/S vssd1 vssd1 vccd1 vccd1 _18795_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15129_ _17897_/Q _15328_/B _15328_/C _12761_/B _15129_/B2 vssd1 vssd1 vccd1 vccd1
+ _15135_/A sky130_fd_sc_hd__a32o_4
XFILLER_217_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09621_ _10315_/S _09621_/B vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__or2_1
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18819_ _19196_/CLK _18819_/D vssd1 vssd1 vccd1 vccd1 _18819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09552_ _09550_/X _09551_/X _09845_/S vssd1 vssd1 vccd1 vccd1 _09553_/B sky130_fd_sc_hd__mux2_1
XFILLER_270_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ _11556_/B _09902_/B vssd1 vssd1 vccd1 vccd1 _09483_/Y sky130_fd_sc_hd__nor2_2
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_86_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17958_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_105_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1307 _15941_/S vssd1 vssd1 vccd1 vccd1 _15947_/S sky130_fd_sc_hd__buf_4
Xfanout1318 _11693_/Y vssd1 vssd1 vccd1 vccd1 _12420_/B1 sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_15_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19602_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout1329 _10004_/A1 vssd1 vssd1 vccd1 vccd1 _10633_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_247_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09819_ _11217_/A _09986_/B _09819_/C vssd1 vssd1 vccd1 vccd1 _09821_/B sky130_fd_sc_hd__and3_1
XFILLER_219_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12830_ _12709_/X _12746_/B _12878_/S vssd1 vssd1 vccd1 vccd1 _12830_/X sky130_fd_sc_hd__mux2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _13185_/A _12761_/B _12761_/C _12761_/D vssd1 vssd1 vccd1 vccd1 _12761_/X
+ sky130_fd_sc_hd__or4_2
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _16470_/A0 _18350_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _18350_/D sky130_fd_sc_hd__mux2_1
XFILLER_203_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11712_ _11712_/A _12271_/A vssd1 vssd1 vccd1 vccd1 _11712_/X sky130_fd_sc_hd__or2_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12688_/X _12691_/X _12943_/S vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__mux2_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15480_ _18118_/Q _15133_/Y _15479_/X _15452_/A vssd1 vssd1 vccd1 vccd1 _15484_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_230_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14431_ _18570_/Q _14450_/B vssd1 vssd1 vccd1 vccd1 _18283_/D sky130_fd_sc_hd__and2_1
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _13740_/B vssd1 vssd1 vccd1 vccd1 _11643_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_230_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17150_ _17261_/A _17150_/B vssd1 vssd1 vccd1 vccd1 _19401_/D sky130_fd_sc_hd__nor2_1
X_14362_ _18214_/Q _17669_/A0 _14382_/S vssd1 vssd1 vccd1 vccd1 _18214_/D sky130_fd_sc_hd__mux2_1
X_11574_ _11327_/S _11573_/X _11572_/X vssd1 vssd1 vccd1 vccd1 _11574_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 core_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
X_16101_ _18753_/Q _16141_/B vssd1 vssd1 vccd1 vccd1 _16101_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput28 core_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10525_ _18126_/Q _10524_/Y _13739_/A vssd1 vssd1 vccd1 vccd1 _12649_/B sky130_fd_sc_hd__mux2_4
X_13313_ _13315_/S _12937_/Y _13413_/B1 vssd1 vssd1 vccd1 vccd1 _13313_/X sky130_fd_sc_hd__a21o_2
Xinput39 core_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17081_ _19374_/Q _17113_/B vssd1 vssd1 vccd1 vccd1 _17081_/X sky130_fd_sc_hd__or2_1
X_14293_ _16611_/A0 _18152_/Q _14305_/S vssd1 vssd1 vccd1 vccd1 _18152_/D sky130_fd_sc_hd__mux2_1
X_16032_ _16020_/Y _16031_/X _16030_/X _16052_/A vssd1 vssd1 vccd1 vccd1 _18729_/D
+ sky130_fd_sc_hd__o211a_1
X_13244_ _19402_/Q _12570_/A _13244_/B1 vssd1 vssd1 vccd1 vccd1 _13244_/X sky130_fd_sc_hd__a21o_1
X_10456_ _10085_/A _10085_/B _09234_/Y _11064_/B1 vssd1 vssd1 vccd1 vccd1 _10456_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_143_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13175_ _15914_/A _12536_/Y _13165_/X _13174_/X _12505_/Y vssd1 vssd1 vccd1 vccd1
+ _13175_/X sky130_fd_sc_hd__a221o_1
XFILLER_272_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10387_ _18465_/Q _18366_/Q _11576_/S vssd1 vssd1 vccd1 vccd1 _10387_/X sky130_fd_sc_hd__mux2_1
XFILLER_272_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12126_ _17836_/Q _12128_/C _12125_/Y vssd1 vssd1 vccd1 vccd1 _17836_/D sky130_fd_sc_hd__o21a_1
X_17983_ _18700_/CLK _17983_/D vssd1 vssd1 vccd1 vccd1 _17983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16934_ _12482_/S _17942_/Q _16933_/X vssd1 vssd1 vccd1 vccd1 _17187_/B sky130_fd_sc_hd__o21a_4
Xfanout1830 _17326_/A vssd1 vssd1 vccd1 vccd1 _14430_/B sky130_fd_sc_hd__buf_4
X_12057_ _17806_/Q _12085_/B vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__or2_1
Xfanout1841 _14181_/A vssd1 vssd1 vccd1 vccd1 _14029_/C1 sky130_fd_sc_hd__buf_4
Xfanout1852 _16904_/A vssd1 vssd1 vccd1 vccd1 _16892_/A sky130_fd_sc_hd__clkbuf_4
Xfanout1863 fanout1870/X vssd1 vssd1 vccd1 vccd1 fanout1863/X sky130_fd_sc_hd__buf_4
X_11008_ _11481_/A _19181_/Q _11395_/C vssd1 vssd1 vccd1 vccd1 _11008_/X sky130_fd_sc_hd__and3_1
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19653_ _19653_/A vssd1 vssd1 vccd1 vccd1 _19653_/X sky130_fd_sc_hd__buf_2
Xfanout1874 _14487_/A vssd1 vssd1 vccd1 vccd1 _16048_/A sky130_fd_sc_hd__buf_8
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1885 fanout1905/X vssd1 vssd1 vccd1 vccd1 _12219_/A sky130_fd_sc_hd__buf_4
X_16865_ _12482_/S _17925_/Q _16864_/X vssd1 vssd1 vccd1 vccd1 _17569_/A sky130_fd_sc_hd__o21a_4
Xfanout1896 _16737_/A vssd1 vssd1 vccd1 vccd1 _16803_/A sky130_fd_sc_hd__clkbuf_4
X_18604_ _19203_/CLK _18604_/D vssd1 vssd1 vccd1 vccd1 _18604_/Q sky130_fd_sc_hd__dfxtp_1
X_15816_ _18608_/Q _16606_/A0 _15833_/S vssd1 vssd1 vccd1 vccd1 _18608_/D sky130_fd_sc_hd__mux2_1
XFILLER_93_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19584_ _19648_/CLK _19584_/D vssd1 vssd1 vccd1 vccd1 _19584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16796_ _19287_/Q _16799_/C _16812_/B1 vssd1 vssd1 vccd1 vccd1 _16796_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18535_ _19148_/CLK _18535_/D vssd1 vssd1 vccd1 vccd1 _18535_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _18591_/Q _15729_/X _15789_/B1 vssd1 vssd1 vccd1 vccd1 _15748_/B sky130_fd_sc_hd__o21ai_1
XFILLER_280_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _12448_/D _12955_/Y _12958_/X _12929_/X vssd1 vssd1 vccd1 vccd1 _12959_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_34_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18466_ _19645_/CLK _18466_/D vssd1 vssd1 vccd1 vccd1 _18466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15678_ _18588_/Q _15704_/C vssd1 vssd1 vccd1 vccd1 _15678_/X sky130_fd_sc_hd__or2_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 input244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_291 _11943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17417_ _18106_/Q _17437_/A2 _17415_/X _17416_/X vssd1 vssd1 vccd1 vccd1 _17417_/X
+ sky130_fd_sc_hd__a22o_1
X_14629_ _17688_/A0 _18436_/Q _14630_/S vssd1 vssd1 vccd1 vccd1 _18436_/D sky130_fd_sc_hd__mux2_1
XFILLER_221_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18397_ _19399_/CLK _18397_/D vssd1 vssd1 vccd1 vccd1 _18397_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17348_ _17360_/A _17348_/B vssd1 vssd1 vccd1 vccd1 _19471_/D sky130_fd_sc_hd__and2_1
XFILLER_159_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17279_ _17277_/Y _17278_/X _16048_/A vssd1 vssd1 vccd1 vccd1 _19443_/D sky130_fd_sc_hd__a21oi_1
XFILLER_228_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19018_ _19640_/CLK _19018_/D vssd1 vssd1 vccd1 vccd1 _19018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08983_ _11428_/A _08982_/X _11501_/B1 vssd1 vssd1 vccd1 vccd1 _08983_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_248_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09604_ _09718_/S _09602_/X _09603_/X _09429_/S vssd1 vssd1 vccd1 vccd1 _09604_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09535_ _09683_/A _09535_/B vssd1 vssd1 vccd1 vccd1 _09535_/X sky130_fd_sc_hd__or2_1
XFILLER_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_133_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19522_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_225_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _09464_/X _09465_/X _10253_/A vssd1 vssd1 vccd1 vccd1 _09466_/X sky130_fd_sc_hd__mux2_1
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09397_ _11046_/S1 _09391_/X _09394_/X _11053_/A vssd1 vssd1 vccd1 vccd1 _09397_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10310_ _17979_/Q _11447_/A2 _11371_/B1 vssd1 vssd1 vccd1 vccd1 _10310_/X sky130_fd_sc_hd__a21o_1
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11290_ _09141_/A _15426_/A _11261_/X vssd1 vssd1 vccd1 vccd1 _12595_/B sky130_fd_sc_hd__o21ai_4
XFILLER_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10241_ _19646_/Q _18935_/Q _10253_/C vssd1 vssd1 vccd1 vccd1 _10241_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10172_ _10253_/A _10170_/X _10171_/X vssd1 vssd1 vccd1 vccd1 _10172_/X sky130_fd_sc_hd__o21a_1
XFILLER_160_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1104 _12589_/X vssd1 vssd1 vccd1 vccd1 _13956_/B1 sky130_fd_sc_hd__buf_6
XFILLER_267_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1115 _12452_/Y vssd1 vssd1 vccd1 vccd1 _13874_/B sky130_fd_sc_hd__buf_4
XFILLER_121_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1126 _12323_/X vssd1 vssd1 vccd1 vccd1 _15661_/B sky130_fd_sc_hd__buf_4
Xfanout1137 _17666_/A0 vssd1 vssd1 vccd1 vccd1 _17699_/A0 sky130_fd_sc_hd__clkbuf_4
X_14980_ _14976_/Y _14979_/X _15010_/B1 vssd1 vssd1 vccd1 vccd1 _14980_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_219_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1148 _09103_/Y vssd1 vssd1 vccd1 vccd1 _11332_/B1 sky130_fd_sc_hd__buf_12
Xfanout1159 _16003_/A2 vssd1 vssd1 vccd1 vccd1 _15977_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13931_ _13931_/A _13931_/B _13931_/C vssd1 vssd1 vccd1 vccd1 _13931_/X sky130_fd_sc_hd__or3_1
XFILLER_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16650_ _19239_/Q _16648_/A _16780_/B1 vssd1 vssd1 vccd1 vccd1 _16651_/B sky130_fd_sc_hd__o21ai_1
XFILLER_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13862_ _11636_/A _13912_/B1 _13912_/A2 _10308_/A _14153_/A vssd1 vssd1 vccd1 vccd1
+ _13862_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_170_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15601_ _15580_/A _15580_/B _15577_/X _15599_/Y _15576_/X vssd1 vssd1 vccd1 vccd1
+ _15620_/B sky130_fd_sc_hd__o311a_1
XFILLER_263_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12813_ _12711_/X _12715_/X _12813_/S vssd1 vssd1 vccd1 vccd1 _12813_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16581_ _16614_/A0 _19185_/Q _16586_/S vssd1 vssd1 vccd1 vccd1 _19185_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13793_ _10604_/Y _13763_/A _13727_/B _12651_/X vssd1 vssd1 vccd1 vccd1 _13794_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_62_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18320_ _19599_/CLK _18320_/D vssd1 vssd1 vccd1 vccd1 _18320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ _15532_/A _15532_/B vssd1 vssd1 vccd1 vccd1 _15536_/B sky130_fd_sc_hd__nor2_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _13315_/S _12746_/B vssd1 vssd1 vccd1 vccd1 _12744_/Y sky130_fd_sc_hd__nor2_1
XFILLER_215_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _19589_/CLK _18251_/D vssd1 vssd1 vccd1 vccd1 _18251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15557_/A _15558_/A vssd1 vssd1 vccd1 vccd1 _15487_/B sky130_fd_sc_hd__nor2_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12675_ _12670_/X _12674_/X _12933_/A vssd1 vssd1 vccd1 vccd1 _12675_/X sky130_fd_sc_hd__mux2_1
XFILLER_231_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17202_ _17202_/A _17202_/B vssd1 vssd1 vccd1 vccd1 _17202_/Y sky130_fd_sc_hd__nand2_2
X_14414_ _17721_/A0 _18265_/Q _14415_/S vssd1 vssd1 vccd1 vccd1 _18265_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11626_ _13962_/A vssd1 vssd1 vccd1 vccd1 _11626_/Y sky130_fd_sc_hd__inv_2
X_18182_ _18613_/CLK _18182_/D vssd1 vssd1 vccd1 vccd1 _18182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15394_ _19437_/Q _15411_/B _17166_/A _15393_/X vssd1 vssd1 vccd1 vccd1 _15394_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ _17157_/A _17567_/A vssd1 vssd1 vccd1 vccd1 _17413_/A sky130_fd_sc_hd__nand2_1
X_14345_ _15039_/A _14345_/B _14345_/C vssd1 vssd1 vccd1 vccd1 _18200_/D sky130_fd_sc_hd__and3_4
XFILLER_128_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11557_ _09048_/A _11556_/X _11219_/B _09987_/A vssd1 vssd1 vccd1 vccd1 _11557_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17064_ _17569_/A _17114_/A2 _17063_/X _17378_/A vssd1 vssd1 vccd1 vccd1 _19365_/D
+ sky130_fd_sc_hd__o211a_1
X_10508_ _19060_/Q _19028_/Q _10656_/S vssd1 vssd1 vccd1 vccd1 _10508_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14276_ _16594_/A0 _18135_/Q _14301_/S vssd1 vssd1 vccd1 vccd1 _18135_/D sky130_fd_sc_hd__mux2_1
X_11488_ _11488_/A _11819_/A vssd1 vssd1 vccd1 vccd1 _11488_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16015_ _18723_/Q _16019_/A2 _16014_/X _14197_/A vssd1 vssd1 vccd1 vccd1 _18723_/D
+ sky130_fd_sc_hd__o211a_1
X_10439_ _10437_/X _10438_/X _10663_/S vssd1 vssd1 vccd1 vccd1 _10439_/X sky130_fd_sc_hd__mux2_1
X_13227_ _13224_/B _13226_/Y _13224_/Y _13227_/C1 vssd1 vssd1 vccd1 vccd1 _13227_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _13150_/X _13157_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _13185_/B sky130_fd_sc_hd__a21oi_1
XFILLER_285_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12109_ _17830_/Q _12112_/C _16149_/A vssd1 vssd1 vccd1 vccd1 _12109_/Y sky130_fd_sc_hd__a21oi_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17966_ _18627_/CLK _17966_/D vssd1 vssd1 vccd1 vccd1 _17966_/Q sky130_fd_sc_hd__dfxtp_1
X_13089_ _13089_/A _13089_/B vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__or2_1
XFILLER_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1660 _11498_/A1 vssd1 vssd1 vccd1 vccd1 _11506_/A1 sky130_fd_sc_hd__clkbuf_8
X_16917_ _18760_/Q _16965_/A2 _16965_/B1 input224/X _16969_/C1 vssd1 vssd1 vccd1 vccd1
+ _16917_/X sky130_fd_sc_hd__a221o_1
XFILLER_266_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1671 _08848_/Y vssd1 vssd1 vccd1 vccd1 _09958_/C1 sky130_fd_sc_hd__buf_12
XFILLER_254_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17897_ _18817_/CLK _17897_/D vssd1 vssd1 vccd1 vccd1 _17897_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1682 _09854_/A vssd1 vssd1 vccd1 vccd1 _11250_/A1 sky130_fd_sc_hd__buf_6
Xfanout1693 _11404_/A1 vssd1 vssd1 vccd1 vccd1 _11389_/A1 sky130_fd_sc_hd__buf_2
XFILLER_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19636_ _19636_/CLK _19636_/D vssd1 vssd1 vccd1 vccd1 _19636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16848_ _08837_/Y _15840_/B _16848_/S vssd1 vssd1 vccd1 vccd1 _16850_/B sky130_fd_sc_hd__mux2_4
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19567_ _19599_/CLK _19567_/D vssd1 vssd1 vccd1 vccd1 _19567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16779_ _16787_/A _16779_/B _16783_/C vssd1 vssd1 vccd1 vccd1 _19280_/D sky130_fd_sc_hd__nor3_1
XFILLER_241_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09320_ input123/X input158/X _09655_/S vssd1 vssd1 vccd1 vccd1 _09320_/X sky130_fd_sc_hd__mux2_8
XFILLER_34_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18518_ _19291_/CLK _18518_/D vssd1 vssd1 vccd1 vccd1 _18518_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_179_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19498_ _19530_/CLK _19498_/D vssd1 vssd1 vccd1 vccd1 _19498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09251_ _09249_/X _09250_/X _10409_/A vssd1 vssd1 vccd1 vccd1 _09251_/X sky130_fd_sc_hd__mux2_1
X_18449_ _19126_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09182_ _10337_/S1 _09181_/X _09180_/X _10338_/A1 vssd1 vssd1 vccd1 vccd1 _09186_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_178_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput207 localMemory_wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput218 localMemory_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input218/X sky130_fd_sc_hd__clkbuf_16
Xinput229 localMemory_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_hd__buf_12
X_08966_ _11497_/A1 _18144_/Q _18790_/Q _08968_/S0 vssd1 vssd1 vccd1 vccd1 _08966_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08897_ _08897_/A _15082_/A vssd1 vssd1 vccd1 vccd1 _08897_/Y sky130_fd_sc_hd__nor2_2
XFILLER_257_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09518_ _11190_/A1 _18210_/Q _09883_/B _18945_/Q _09723_/S vssd1 vssd1 vccd1 vccd1
+ _09518_/X sky130_fd_sc_hd__o221a_1
X_10790_ _10781_/Y _10788_/Y _10789_/X _10775_/X vssd1 vssd1 vccd1 vccd1 _10790_/X
+ sky130_fd_sc_hd__o2bb2a_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _10263_/A1 _19561_/Q _10249_/S _19593_/Q _10266_/S1 vssd1 vssd1 vccd1 vccd1
+ _09449_/X sky130_fd_sc_hd__o221a_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12460_ _12460_/A _13289_/A vssd1 vssd1 vccd1 vccd1 _12460_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _11411_/A _11823_/A vssd1 vssd1 vccd1 vccd1 _11411_/Y sky130_fd_sc_hd__nor2_1
X_12391_ _12430_/A _12391_/B vssd1 vssd1 vccd1 vccd1 _12391_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11342_ _11355_/A1 _11341_/X _11623_/A1 vssd1 vssd1 vccd1 vccd1 _11342_/X sky130_fd_sc_hd__a21o_1
X_14130_ _16547_/A0 _18069_/Q _14140_/S vssd1 vssd1 vccd1 vccd1 _18069_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18445_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14061_ _17678_/A0 _18003_/Q _14073_/S vssd1 vssd1 vccd1 vccd1 _18003_/D sky130_fd_sc_hd__mux2_1
X_11273_ _10745_/S _11270_/X _11272_/X vssd1 vssd1 vccd1 vccd1 _11273_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_141_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13012_ _17828_/Q _13944_/B vssd1 vssd1 vccd1 vccd1 _13012_/X sky130_fd_sc_hd__or2_1
X_10224_ _19647_/Q _18936_/Q _10224_/S vssd1 vssd1 vccd1 vccd1 _10224_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17820_ _19492_/CLK _17820_/D vssd1 vssd1 vccd1 vccd1 _17820_/Q sky130_fd_sc_hd__dfxtp_4
X_10155_ _11518_/B2 _10089_/B _10154_/Y _11055_/B2 vssd1 vssd1 vccd1 vccd1 _13917_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_67_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17751_ _18651_/Q vssd1 vssd1 vccd1 vccd1 _18651_/D sky130_fd_sc_hd__clkbuf_2
X_10086_ _10086_/A _10309_/B vssd1 vssd1 vccd1 vccd1 _10086_/Y sky130_fd_sc_hd__nor2_1
X_14963_ _14992_/A1 _13831_/Y _14973_/B1 _18653_/Q _14973_/C1 vssd1 vssd1 vccd1 vccd1
+ _14963_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16702_ _19253_/Q _16708_/D _16701_/Y _16964_/A vssd1 vssd1 vccd1 vccd1 _19253_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_208_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13914_ _12442_/D _12835_/B _14155_/B _12656_/A _13913_/X vssd1 vssd1 vccd1 vccd1
+ _13914_/X sky130_fd_sc_hd__o221a_1
X_17682_ _17682_/A0 _19609_/Q _17690_/S vssd1 vssd1 vccd1 vccd1 _19609_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14894_ _14854_/X _14893_/X _14726_/X vssd1 vssd1 vccd1 vccd1 _16078_/C sky130_fd_sc_hd__a21oi_2
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19421_ _19453_/CLK _19421_/D vssd1 vssd1 vccd1 vccd1 _19421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16633_ _17724_/A _19233_/Q _19232_/Q vssd1 vssd1 vccd1 vccd1 _16677_/A sky130_fd_sc_hd__and3_2
X_13845_ _19260_/Q _13943_/A2 _13943_/B1 _19292_/Q vssd1 vssd1 vccd1 vccd1 _13845_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_223_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19352_ _19483_/CLK _19352_/D vssd1 vssd1 vccd1 vccd1 _19352_/Q sky130_fd_sc_hd__dfxtp_1
X_16564_ _17697_/A0 _19168_/Q _16586_/S vssd1 vssd1 vccd1 vccd1 _19168_/D sky130_fd_sc_hd__mux2_1
X_13776_ _17849_/Q _13844_/A2 _13844_/B1 _17881_/Q vssd1 vssd1 vccd1 vccd1 _13776_/X
+ sky130_fd_sc_hd__a22o_1
X_10988_ _10988_/A _10988_/B vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18303_ _19453_/CLK _18303_/D vssd1 vssd1 vccd1 vccd1 _18303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15515_ _15789_/A1 _15511_/Y _15537_/B1 vssd1 vssd1 vccd1 vccd1 _15515_/Y sky130_fd_sc_hd__a21oi_1
X_19283_ _19295_/CLK _19283_/D vssd1 vssd1 vccd1 vccd1 _19283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12727_ _12722_/X _12726_/Y _12933_/A vssd1 vssd1 vccd1 vccd1 _12727_/X sky130_fd_sc_hd__mux2_1
X_16495_ _16594_/A0 _19101_/Q _16515_/S vssd1 vssd1 vccd1 vccd1 _19101_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18234_ _19225_/CLK _18234_/D vssd1 vssd1 vccd1 vccd1 _18234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15446_ _15498_/S _15445_/Y _15440_/Y _17166_/A vssd1 vssd1 vccd1 vccd1 _15446_/X
+ sky130_fd_sc_hd__a211o_1
X_12658_ _10307_/A _12658_/B vssd1 vssd1 vccd1 vccd1 _12658_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11609_ _18338_/Q _17789_/Q _11609_/S vssd1 vssd1 vccd1 vccd1 _11609_/X sky130_fd_sc_hd__mux2_1
X_18165_ _18875_/CLK _18165_/D vssd1 vssd1 vccd1 vccd1 _18165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15377_ _19468_/Q _15376_/X _15498_/S vssd1 vssd1 vccd1 vccd1 _15377_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12589_ _12754_/B _12455_/A _12587_/B vssd1 vssd1 vccd1 vccd1 _12589_/X sky130_fd_sc_hd__o21a_1
XFILLER_239_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17116_ _17214_/B _17116_/A2 _17115_/X _17354_/A vssd1 vssd1 vccd1 vccd1 _19391_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14328_ _18185_/Q _16314_/A0 _14339_/S vssd1 vssd1 vccd1 vccd1 _18185_/D sky130_fd_sc_hd__mux2_1
X_18096_ _18761_/CLK _18096_/D vssd1 vssd1 vccd1 vccd1 _18096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17047_ _17051_/A _17047_/B vssd1 vssd1 vccd1 vccd1 _17381_/C sky130_fd_sc_hd__or2_4
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14259_ _18301_/Q _14261_/A2 _14258_/X _14451_/B vssd1 vssd1 vccd1 vccd1 _18127_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 _16425_/S vssd1 vssd1 vccd1 vccd1 _16420_/S sky130_fd_sc_hd__buf_12
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout919 _16260_/Y vssd1 vssd1 vccd1 vccd1 _16278_/S sky130_fd_sc_hd__buf_8
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08820_ _19427_/Q vssd1 vssd1 vccd1 vccd1 _08820_/Y sky130_fd_sc_hd__inv_2
XFILLER_285_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18998_ _19596_/CLK _18998_/D vssd1 vssd1 vccd1 vccd1 _18998_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _17951_/CLK _17949_/D vssd1 vssd1 vccd1 vccd1 _17949_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1490 _10721_/S vssd1 vssd1 vccd1 vccd1 _10370_/S sky130_fd_sc_hd__buf_6
XFILLER_241_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19619_ _19619_/CLK _19619_/D vssd1 vssd1 vccd1 vccd1 _19619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09303_ _18635_/Q _18057_/Q _09306_/S vssd1 vssd1 vccd1 vccd1 _09303_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _11218_/A _09902_/C vssd1 vssd1 vccd1 vccd1 _09234_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09165_ _11469_/A1 _17768_/Q _09179_/B _18317_/Q _10338_/A1 vssd1 vssd1 vccd1 vccd1
+ _09165_/X sky130_fd_sc_hd__o221a_1
XFILLER_210_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ _11251_/S _12442_/B vssd1 vssd1 vccd1 vccd1 _09096_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09998_ _11157_/A1 _19554_/Q _11154_/S _19586_/Q _11569_/S1 vssd1 vssd1 vccd1 vccd1
+ _09998_/X sky130_fd_sc_hd__o221a_1
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ _10275_/S _14074_/B vssd1 vssd1 vccd1 vccd1 _08956_/B sky130_fd_sc_hd__xnor2_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11960_ _18506_/Q _11720_/X _11910_/X _11706_/X vssd1 vssd1 vccd1 vccd1 _11960_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10911_ _17971_/Q _11216_/A2 _11216_/B1 vssd1 vssd1 vccd1 vccd1 _10912_/B sky130_fd_sc_hd__a21oi_1
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11891_ _10271_/B _11864_/B _11952_/A2 vssd1 vssd1 vccd1 vccd1 _11894_/B sky130_fd_sc_hd__o21ai_2
XFILLER_244_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13630_ _19413_/Q _13654_/A2 _13654_/B1 vssd1 vssd1 vccd1 vccd1 _13630_/X sky130_fd_sc_hd__a21o_1
XFILLER_204_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10842_ _10850_/A1 _18224_/Q _11581_/S _18959_/Q _10918_/C1 vssd1 vssd1 vccd1 vccd1
+ _10842_/X sky130_fd_sc_hd__o221a_1
XFILLER_13_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13561_ _14012_/B vssd1 vssd1 vccd1 vccd1 _13561_/Y sky130_fd_sc_hd__inv_2
X_10773_ _18154_/Q _11482_/A2 _10772_/X _11578_/S vssd1 vssd1 vccd1 vccd1 _10773_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_200_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15300_ _19465_/Q _15299_/Y _15498_/S vssd1 vssd1 vccd1 vccd1 _15300_/X sky130_fd_sc_hd__mux2_1
XFILLER_212_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ _12563_/A _12512_/B vssd1 vssd1 vccd1 vccd1 _12768_/A sky130_fd_sc_hd__nand2b_4
XFILLER_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16280_ _16611_/A0 _18894_/Q _16292_/S vssd1 vssd1 vccd1 vccd1 _18894_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13492_ _15478_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _13507_/B sky130_fd_sc_hd__or2_1
XFILLER_200_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15231_ _19461_/Q _19395_/Q _15204_/B vssd1 vssd1 vccd1 vccd1 _15231_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12443_ _12443_/A _12443_/B _12443_/C _12443_/D vssd1 vssd1 vccd1 vccd1 _12445_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_138_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15162_ _08820_/Y _15416_/A _15731_/B1 _15161_/Y _17219_/A vssd1 vssd1 vccd1 vccd1
+ _15163_/B sky130_fd_sc_hd__a221o_1
X_12374_ _17899_/Q _12421_/A _12373_/Y _12428_/C1 vssd1 vssd1 vccd1 vccd1 _17899_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14113_ _17663_/A0 _18052_/Q _14131_/S vssd1 vssd1 vccd1 vccd1 _18052_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11325_ _18857_/Q _18889_/Q _11325_/S vssd1 vssd1 vccd1 vccd1 _11325_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15093_ _15093_/A _15093_/B _15093_/C _15093_/D vssd1 vssd1 vccd1 vccd1 _17591_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_114_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18921_ _19632_/CLK _18921_/D vssd1 vssd1 vccd1 vccd1 _18921_/Q sky130_fd_sc_hd__dfxtp_1
X_14044_ _17694_/A0 _17986_/Q _14064_/S vssd1 vssd1 vccd1 vccd1 _17986_/D sky130_fd_sc_hd__mux2_1
X_11256_ _11254_/X _11255_/X _11332_/B1 vssd1 vssd1 vccd1 vccd1 _11256_/X sky130_fd_sc_hd__a21o_2
XFILLER_192_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10207_ _10354_/A1 _18233_/Q _10206_/S _18968_/Q _10205_/S vssd1 vssd1 vccd1 vccd1
+ _10207_/X sky130_fd_sc_hd__o221a_1
XFILLER_192_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18852_ _19627_/CLK _18852_/D vssd1 vssd1 vccd1 vccd1 _18852_/Q sky130_fd_sc_hd__dfxtp_1
X_11187_ _09723_/S _11186_/X _11515_/B1 vssd1 vssd1 vccd1 vccd1 _11187_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_279_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10138_ _19065_/Q _19033_/Q _10224_/S vssd1 vssd1 vccd1 vccd1 _10138_/X sky130_fd_sc_hd__mux2_1
X_17803_ _17930_/CLK _17803_/D vssd1 vssd1 vccd1 vccd1 _17803_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_269_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18783_ _19138_/CLK _18783_/D vssd1 vssd1 vccd1 vccd1 _18783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ _18713_/Q _16003_/A2 _15994_/X _14203_/A vssd1 vssd1 vccd1 vccd1 _18713_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17734_ _18634_/Q vssd1 vssd1 vccd1 vccd1 _18634_/D sky130_fd_sc_hd__clkbuf_2
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14946_ _15006_/A1 _14945_/X _15006_/B1 vssd1 vssd1 vccd1 vccd1 _14946_/Y sky130_fd_sc_hd__o21ai_2
X_10069_ _11731_/B _10068_/B _11734_/B vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__a21o_1
XFILLER_75_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17665_ _17665_/A0 _19592_/Q _17687_/S vssd1 vssd1 vccd1 vccd1 _19592_/D sky130_fd_sc_hd__mux2_1
X_14877_ _14877_/A vssd1 vssd1 vccd1 vccd1 _14877_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19404_ _19464_/CLK _19404_/D vssd1 vssd1 vccd1 vccd1 _19404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16616_ _17683_/A0 _19219_/Q _16618_/S vssd1 vssd1 vccd1 vccd1 _19219_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13828_ _19387_/Q _13884_/A2 _13826_/X _13827_/X _13884_/C1 vssd1 vssd1 vccd1 vccd1
+ _13828_/X sky130_fd_sc_hd__o221a_4
X_17596_ _19539_/Q _17622_/A2 _17591_/X _17172_/B _17595_/X vssd1 vssd1 vccd1 vccd1
+ _19539_/D sky130_fd_sc_hd__o221a_1
XFILLER_91_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19335_ _19464_/CLK _19335_/D vssd1 vssd1 vccd1 vccd1 _19335_/Q sky130_fd_sc_hd__dfxtp_1
X_16547_ _16547_/A0 _19152_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _19152_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13759_ _13758_/B _13757_/X _13758_/Y _13930_/B1 _13931_/A vssd1 vssd1 vccd1 vccd1
+ _13759_/X sky130_fd_sc_hd__a221o_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19266_ _19268_/CLK _19266_/D vssd1 vssd1 vccd1 vccd1 _19266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16478_ _17677_/A0 _19085_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _19085_/D sky130_fd_sc_hd__mux2_1
X_18217_ _19612_/CLK _18217_/D vssd1 vssd1 vccd1 vccd1 _18217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15429_ _09494_/A _15429_/A2 _15484_/A vssd1 vssd1 vccd1 vccd1 _15432_/B sky130_fd_sc_hd__o21a_2
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19197_ _19197_/CLK _19197_/D vssd1 vssd1 vccd1 vccd1 _19197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18148_ _19025_/CLK _18148_/D vssd1 vssd1 vccd1 vccd1 _18148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18079_ _19163_/CLK _18079_/D vssd1 vssd1 vccd1 vccd1 _18079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09921_ _10262_/A1 _18205_/Q _09925_/S _18940_/Q _10266_/S1 vssd1 vssd1 vccd1 vccd1
+ _09921_/X sky130_fd_sc_hd__o221a_1
XFILLER_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout705 _12543_/X vssd1 vssd1 vccd1 vccd1 _13846_/B sky130_fd_sc_hd__buf_6
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout716 _12541_/Y vssd1 vssd1 vccd1 vccd1 _12919_/A2 sky130_fd_sc_hd__buf_4
Xfanout727 _12495_/Y vssd1 vssd1 vccd1 vccd1 _13164_/A2 sky130_fd_sc_hd__buf_2
X_09852_ _18309_/Q _17760_/Q _11147_/S vssd1 vssd1 vccd1 vccd1 _09852_/X sky130_fd_sc_hd__mux2_1
XFILLER_258_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout738 _16507_/A0 vssd1 vssd1 vccd1 vccd1 _16540_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_112_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout749 _13046_/A1 vssd1 vssd1 vccd1 vccd1 _13354_/A sky130_fd_sc_hd__buf_4
XFILLER_259_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _10036_/S _09782_/X _09781_/X vssd1 vssd1 vccd1 vccd1 _09783_/X sky130_fd_sc_hd__o21a_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_109 _11737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09217_ _09215_/X _09216_/X _10205_/S vssd1 vssd1 vccd1 vccd1 _09217_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09148_ _11218_/A _09819_/C vssd1 vssd1 vccd1 vccd1 _09148_/X sky130_fd_sc_hd__or2_1
XFILLER_135_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ _12443_/A _09080_/B _09080_/C vssd1 vssd1 vccd1 vccd1 _09079_/Y sky130_fd_sc_hd__nor3_4
XFILLER_163_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11110_ _11355_/A1 _11109_/X _11608_/C1 vssd1 vssd1 vccd1 vccd1 _11110_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_146_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_3__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_3__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ _12035_/B _12089_/Y _14487_/A vssd1 vssd1 vccd1 vccd1 _17822_/D sky130_fd_sc_hd__a21o_1
XFILLER_104_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11041_ _11498_/A1 _18151_/Q _18797_/Q _09966_/S vssd1 vssd1 vccd1 vccd1 _11041_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _17801_/Q _14799_/X _14993_/S vssd1 vssd1 vccd1 vccd1 _14800_/X sky130_fd_sc_hd__mux2_1
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _15780_/A _15780_/B vssd1 vssd1 vccd1 vccd1 _15780_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_58_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12992_ _12992_/A vssd1 vssd1 vccd1 vccd1 _12992_/Y sky130_fd_sc_hd__inv_2
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _18474_/Q _14720_/A _14730_/Y _17159_/A vssd1 vssd1 vccd1 vccd1 _18474_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_18_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11943_ _11944_/A1 _11872_/B _11959_/A2 input230/X vssd1 vssd1 vccd1 vccd1 _11943_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _11683_/B _17475_/A2 _17475_/B1 _17802_/Q _15116_/B vssd1 vssd1 vccd1 vccd1
+ _17450_/X sky130_fd_sc_hd__a221o_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _17721_/A0 _18468_/Q _14663_/S vssd1 vssd1 vccd1 vccd1 _18468_/D sky130_fd_sc_hd__mux2_1
XFILLER_229_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11874_ _12842_/A _14141_/B vssd1 vssd1 vccd1 vccd1 _11901_/B sky130_fd_sc_hd__nand2_8
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _17666_/A0 _19010_/Q _16424_/S vssd1 vssd1 vccd1 vccd1 _19010_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _17940_/Q _13742_/A2 _13612_/X _14177_/A vssd1 vssd1 vccd1 vccd1 _17940_/D
+ sky130_fd_sc_hd__o211a_1
X_17381_ _17555_/B _17381_/B _17381_/C vssd1 vssd1 vccd1 vccd1 _17382_/B sky130_fd_sc_hd__nor3_4
XFILLER_38_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10825_ _08874_/D _10824_/X _11608_/C1 vssd1 vssd1 vccd1 vccd1 _10825_/X sky130_fd_sc_hd__a21o_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14593_ _11706_/C _11818_/B _08884_/X vssd1 vssd1 vccd1 vccd1 _14593_/X sky130_fd_sc_hd__a21o_1
XFILLER_158_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19120_ _19649_/CLK _19120_/D vssd1 vssd1 vccd1 vccd1 _19120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16332_ _18944_/Q _17664_/A0 _16352_/S vssd1 vssd1 vccd1 vccd1 _18944_/D sky130_fd_sc_hd__mux2_1
X_13544_ _13904_/A _13544_/B vssd1 vssd1 vccd1 vccd1 _13544_/Y sky130_fd_sc_hd__nand2_1
X_10756_ _09034_/B _09572_/X _09326_/A vssd1 vssd1 vccd1 vccd1 _10757_/B sky130_fd_sc_hd__a21oi_1
XFILLER_200_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19051_ _19622_/CLK _19051_/D vssd1 vssd1 vccd1 vccd1 _19051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16263_ _16594_/A0 _18877_/Q _16288_/S vssd1 vssd1 vccd1 vccd1 _18877_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13475_ _13545_/A _13475_/B vssd1 vssd1 vccd1 vccd1 _13475_/Y sky130_fd_sc_hd__nand2_1
XFILLER_200_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10687_ _19057_/Q _19025_/Q _10687_/S vssd1 vssd1 vccd1 vccd1 _10687_/X sky130_fd_sc_hd__mux2_1
X_18002_ _19636_/CLK _18002_/D vssd1 vssd1 vccd1 vccd1 _18002_/Q sky130_fd_sc_hd__dfxtp_1
X_15214_ _15214_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _15214_/X sky130_fd_sc_hd__and2_1
X_12426_ _12429_/A1 _12432_/A2 _09569_/X _12429_/B1 _18402_/Q vssd1 vssd1 vccd1 vccd1
+ _12427_/B sky130_fd_sc_hd__o32ai_4
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16194_ _16359_/A _16194_/B vssd1 vssd1 vccd1 vccd1 _16194_/X sky130_fd_sc_hd__or2_4
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput308 _11756_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[12] sky130_fd_sc_hd__buf_4
X_15145_ _17157_/A _15145_/B _15145_/C vssd1 vssd1 vccd1 vccd1 _15145_/X sky130_fd_sc_hd__or3_1
X_12357_ _11695_/B _09991_/A _09477_/X _12432_/B1 _18379_/Q vssd1 vssd1 vccd1 vccd1
+ _12358_/B sky130_fd_sc_hd__o32ai_4
XFILLER_114_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput319 _11766_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[22] sky130_fd_sc_hd__buf_4
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11308_ _18421_/Q _11300_/B _11307_/X _10784_/S vssd1 vssd1 vccd1 vccd1 _11308_/X
+ sky130_fd_sc_hd__o211a_1
X_15076_ _18560_/Q _16488_/A0 _15076_/S vssd1 vssd1 vccd1 vccd1 _18560_/D sky130_fd_sc_hd__mux2_1
X_12288_ _18096_/Q _12305_/A2 _12305_/B1 _18519_/Q vssd1 vssd1 vccd1 vccd1 _12457_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_206_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18904_ _19193_/CLK _18904_/D vssd1 vssd1 vccd1 vccd1 _18904_/Q sky130_fd_sc_hd__dfxtp_1
X_14027_ _17978_/Q _14027_/A2 _14026_/Y _14029_/C1 vssd1 vssd1 vccd1 vccd1 _17978_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11239_ _19633_/Q _18922_/Q _11247_/S vssd1 vssd1 vccd1 vccd1 _11239_/X sky130_fd_sc_hd__mux2_1
XFILLER_267_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18835_ _19641_/CLK _18835_/D vssd1 vssd1 vccd1 vccd1 _18835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18766_ _19076_/CLK _18766_/D vssd1 vssd1 vccd1 vccd1 _18766_/Q sky130_fd_sc_hd__dfxtp_1
X_15978_ _18704_/Q _15953_/B _16004_/B1 _18753_/Q _16018_/C1 vssd1 vssd1 vccd1 vccd1
+ _15978_/X sky130_fd_sc_hd__a221o_1
XFILLER_209_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14929_ _14925_/Y _14928_/X _14950_/B1 vssd1 vssd1 vccd1 vccd1 _14929_/Y sky130_fd_sc_hd__a21oi_4
X_17717_ _17717_/A0 _19643_/Q _17718_/S vssd1 vssd1 vccd1 vccd1 _19643_/D sky130_fd_sc_hd__mux2_1
XFILLER_282_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18697_ _19304_/CLK _18697_/D vssd1 vssd1 vccd1 vccd1 _18697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17648_ _17681_/A0 _19576_/Q _17648_/S vssd1 vssd1 vccd1 vccd1 _19576_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17579_ _17579_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17579_/X sky130_fd_sc_hd__or2_1
XFILLER_251_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19318_ _19319_/CLK _19318_/D vssd1 vssd1 vccd1 vccd1 _19318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19249_ _19268_/CLK _19249_/D vssd1 vssd1 vccd1 vccd1 _19249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09002_ input113/X input148/X _09651_/S vssd1 vssd1 vccd1 vccd1 _09002_/X sky130_fd_sc_hd__mux2_8
XFILLER_192_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_158_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19531_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09904_ _09245_/A _09903_/X _09900_/Y vssd1 vssd1 vccd1 vccd1 _09904_/Y sky130_fd_sc_hd__a21oi_1
Xfanout502 _11959_/B2 vssd1 vssd1 vccd1 vccd1 _11944_/A1 sky130_fd_sc_hd__buf_4
Xfanout513 _17389_/X vssd1 vssd1 vccd1 vccd1 _17499_/A2 sky130_fd_sc_hd__buf_6
XFILLER_263_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout524 _15127_/Y vssd1 vssd1 vccd1 vccd1 _15447_/B sky130_fd_sc_hd__buf_6
Xfanout535 fanout536/X vssd1 vssd1 vccd1 vccd1 _17124_/B sky130_fd_sc_hd__buf_2
XFILLER_258_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout546 _17389_/B1 vssd1 vssd1 vccd1 vccd1 _17382_/A sky130_fd_sc_hd__buf_4
XFILLER_274_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout557 _15787_/A vssd1 vssd1 vccd1 vccd1 _15744_/A sky130_fd_sc_hd__buf_4
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09835_ _19037_/Q _19005_/Q _11147_/S vssd1 vssd1 vccd1 vccd1 _09835_/X sky130_fd_sc_hd__mux2_1
Xfanout568 _15623_/A vssd1 vssd1 vccd1 vccd1 _15369_/A sky130_fd_sc_hd__buf_8
Xfanout579 _12421_/A vssd1 vssd1 vccd1 vccd1 _12408_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_281_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09766_ _11084_/S _09765_/X _11570_/B1 vssd1 vssd1 vccd1 vccd1 _09766_/X sky130_fd_sc_hd__o21a_1
XFILLER_273_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _11252_/S _09697_/B vssd1 vssd1 vccd1 vccd1 _09697_/Y sky130_fd_sc_hd__nand2_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10610_ _19641_/Q _18930_/Q _10619_/S vssd1 vssd1 vccd1 vccd1 _10610_/X sky130_fd_sc_hd__mux2_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11590_ _10399_/A _11571_/Y _11589_/X vssd1 vssd1 vccd1 vccd1 _11590_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_195_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _18260_/Q _18835_/Q _10619_/S vssd1 vssd1 vccd1 vccd1 _10541_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13260_ _13260_/A _13260_/B vssd1 vssd1 vccd1 vccd1 _13260_/Y sky130_fd_sc_hd__nand2_1
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10472_ _10462_/X _10465_/X _10468_/X _10471_/X _11583_/A _11588_/B1 vssd1 vssd1
+ vccd1 vccd1 _10473_/B sky130_fd_sc_hd__mux4_2
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12211_ _16811_/A _12216_/C vssd1 vssd1 vccd1 vccd1 _12211_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13191_ _11751_/A _13483_/B _13190_/Y vssd1 vssd1 vccd1 vccd1 _13191_/X sky130_fd_sc_hd__a21o_1
XFILLER_157_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _17842_/Q _12144_/C _12141_/Y vssd1 vssd1 vccd1 vccd1 _17842_/D sky130_fd_sc_hd__o21a_1
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16950_ _16970_/A1 _17946_/Q _16949_/X vssd1 vssd1 vccd1 vccd1 _17199_/B sky130_fd_sc_hd__o21a_4
XFILLER_173_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12073_ _17814_/Q _12073_/B vssd1 vssd1 vccd1 vccd1 _12073_/X sky130_fd_sc_hd__or2_1
XFILLER_2_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15901_ _18676_/Q _15910_/A2 _15900_/X _15904_/C1 vssd1 vssd1 vccd1 vccd1 _18676_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_249_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11024_ _11024_/A1 _11022_/X _11023_/X vssd1 vssd1 vccd1 vccd1 _11845_/A sky130_fd_sc_hd__o21ai_4
X_16881_ _18751_/Q _16893_/A2 _16893_/B1 input246/X _12483_/A vssd1 vssd1 vccd1 vccd1
+ _16881_/X sky130_fd_sc_hd__a221o_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15832_ _18624_/Q _15832_/A1 _15832_/S vssd1 vssd1 vccd1 vccd1 _18624_/D sky130_fd_sc_hd__mux2_1
X_18620_ _19644_/CLK _18620_/D vssd1 vssd1 vccd1 vccd1 _18620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _18131_/Q _15763_/A2 _15762_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _15765_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_18_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18551_ _19600_/CLK _18551_/D vssd1 vssd1 vccd1 vccd1 _18551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12975_ _15869_/A _12506_/X _12964_/X _12974_/X _12510_/X vssd1 vssd1 vccd1 vccd1
+ _12977_/A sky130_fd_sc_hd__o221a_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _14714_/A _14714_/B vssd1 vssd1 vccd1 vccd1 _14714_/Y sky130_fd_sc_hd__nand2_1
X_17502_ _18123_/Q _17545_/C1 _17500_/X _17501_/X vssd1 vssd1 vccd1 vccd1 _17502_/X
+ sky130_fd_sc_hd__a22o_1
X_18482_ _18517_/CLK _18482_/D vssd1 vssd1 vccd1 vccd1 _18482_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _11926_/A1 _11939_/A1 _11865_/B _11935_/B1 input243/X vssd1 vssd1 vccd1 vccd1
+ _11926_/X sky130_fd_sc_hd__a32o_4
XFILLER_206_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15694_ _19482_/Q _19416_/Q vssd1 vssd1 vccd1 vccd1 _15695_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_440 _13157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_451 _13808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_462 _18384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17433_ _17433_/A _17462_/B vssd1 vssd1 vccd1 vccd1 _17433_/Y sky130_fd_sc_hd__nand2_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _17704_/A0 _18451_/Q _14663_/S vssd1 vssd1 vccd1 vccd1 _18451_/D sky130_fd_sc_hd__mux2_1
XFILLER_205_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_473 input219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11857_ _11909_/A _11857_/B vssd1 vssd1 vccd1 vccd1 _11857_/X sky130_fd_sc_hd__and2_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_484 _11924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_495 _11955_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17364_ _17368_/A _17364_/B vssd1 vssd1 vccd1 vccd1 _19479_/D sky130_fd_sc_hd__and2_1
X_10808_ _11357_/S1 _10797_/X _10807_/X _11621_/C1 vssd1 vssd1 vccd1 vccd1 _10808_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14576_ _14576_/A _14576_/B vssd1 vssd1 vccd1 vccd1 _18396_/D sky130_fd_sc_hd__or2_1
X_11788_ _11816_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11846_/B sky130_fd_sc_hd__nor2_8
X_19103_ _19201_/CLK _19103_/D vssd1 vssd1 vccd1 vccd1 _19103_/Q sky130_fd_sc_hd__dfxtp_1
X_16315_ _17713_/A0 _18928_/Q _16320_/S vssd1 vssd1 vccd1 vccd1 _18928_/D sky130_fd_sc_hd__mux2_1
X_13527_ _13517_/Y _13526_/Y _13527_/B1 _13516_/X vssd1 vssd1 vccd1 vccd1 _13527_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17295_ _19449_/Q _17307_/B vssd1 vssd1 vccd1 vccd1 _17295_/Y sky130_fd_sc_hd__nand2_1
X_10739_ _11277_/A1 _18155_/Q _18801_/Q _10744_/S vssd1 vssd1 vccd1 vccd1 _10739_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19034_ _19118_/CLK _19034_/D vssd1 vssd1 vccd1 vccd1 _19034_/Q sky130_fd_sc_hd__dfxtp_1
X_16246_ _16610_/A0 _18861_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _18861_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13458_ _13527_/B1 _13447_/X _13449_/Y _13457_/Y vssd1 vssd1 vccd1 vccd1 _14006_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12409_ _11695_/B _12409_/A2 _09008_/X _12432_/B1 _18396_/Q vssd1 vssd1 vccd1 vccd1
+ _12409_/X sky130_fd_sc_hd__o32a_1
X_16177_ _16607_/A0 _18794_/Q _16189_/S vssd1 vssd1 vccd1 vccd1 _18794_/D sky130_fd_sc_hd__mux2_1
X_13389_ _13086_/X _13090_/Y _13414_/A vssd1 vssd1 vccd1 vccd1 _13389_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15128_ _15108_/A _15108_/B _15108_/X _15109_/X vssd1 vssd1 vccd1 vccd1 _15137_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_217_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15059_ _18543_/Q _17670_/A0 _15078_/S vssd1 vssd1 vccd1 vccd1 _18543_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09620_ _09618_/X _09619_/X _10706_/S vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__mux2_1
X_18818_ _18880_/CLK _18818_/D vssd1 vssd1 vccd1 vccd1 _18818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09551_ _19624_/Q _18913_/Q _09925_/S vssd1 vssd1 vccd1 vccd1 _09551_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18749_ _18749_/CLK _18749_/D vssd1 vssd1 vccd1 vccd1 _18749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09482_ _18387_/Q _09656_/B1 _09331_/A _09481_/Y vssd1 vssd1 vccd1 vccd1 _09489_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1308 _15881_/B vssd1 vssd1 vccd1 vccd1 _15941_/S sky130_fd_sc_hd__buf_4
XFILLER_266_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1319 _09457_/Y vssd1 vssd1 vccd1 vccd1 _11482_/A2 sky130_fd_sc_hd__buf_12
XFILLER_275_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09818_ _13263_/A _09818_/B vssd1 vssd1 vccd1 vccd1 _11734_/B sky130_fd_sc_hd__nor2_4
XFILLER_275_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_55_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19647_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_274_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09749_ _09747_/X _09748_/X _11568_/A vssd1 vssd1 vccd1 vccd1 _09749_/X sky130_fd_sc_hd__mux2_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12665_/X _12758_/X _12759_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _12761_/D
+ sky130_fd_sc_hd__a31oi_2
XFILLER_199_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11711_/A _11711_/B vssd1 vssd1 vccd1 vccd1 _12271_/A sky130_fd_sc_hd__nand2_4
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12691_ _12689_/X _12690_/X _12796_/S vssd1 vssd1 vccd1 vccd1 _12691_/X sky130_fd_sc_hd__mux2_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _18569_/Q _14430_/B vssd1 vssd1 vccd1 vccd1 _18282_/D sky130_fd_sc_hd__and2_1
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11642_ _13727_/A _11642_/B vssd1 vssd1 vccd1 vccd1 _13740_/B sky130_fd_sc_hd__xnor2_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14361_ _18213_/Q _16535_/A0 _14382_/S vssd1 vssd1 vccd1 vccd1 _18213_/D sky130_fd_sc_hd__mux2_1
X_11573_ _18874_/Q _18906_/Q _11576_/S vssd1 vssd1 vccd1 vccd1 _11573_/X sky130_fd_sc_hd__mux2_1
X_16100_ _16142_/A1 _16099_/Y _16149_/A vssd1 vssd1 vccd1 vccd1 _18752_/D sky130_fd_sc_hd__a21oi_1
XFILLER_156_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 core_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
X_13312_ _13312_/A _14144_/B vssd1 vssd1 vccd1 vccd1 _13312_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17080_ _17585_/A _17114_/A2 _17079_/X _17346_/A vssd1 vssd1 vccd1 vccd1 _19373_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10524_ _13743_/A vssd1 vssd1 vccd1 vccd1 _10524_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 core_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_2
X_14292_ _16610_/A0 _18151_/Q _14304_/S vssd1 vssd1 vccd1 vccd1 _18151_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16031_ _18736_/Q _18728_/Q _16034_/S vssd1 vssd1 vccd1 vccd1 _16031_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13243_ _19500_/Q _13064_/B _13243_/B1 _13242_/X vssd1 vssd1 vccd1 vccd1 _13243_/X
+ sky130_fd_sc_hd__o211a_1
X_10455_ _11639_/A vssd1 vssd1 vccd1 vccd1 _13794_/A sky130_fd_sc_hd__clkinv_4
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13174_ _13174_/A _13174_/B _13174_/C vssd1 vssd1 vccd1 vccd1 _13174_/X sky130_fd_sc_hd__or3_4
XFILLER_123_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10386_ _19644_/Q _18933_/Q _11576_/S vssd1 vssd1 vccd1 vccd1 _10386_/X sky130_fd_sc_hd__mux2_1
XFILLER_269_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12125_ _17836_/Q _12128_/C _12219_/A vssd1 vssd1 vccd1 vccd1 _12125_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17982_ _17982_/CLK _17982_/D vssd1 vssd1 vccd1 vccd1 _17982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1820 fanout1870/X vssd1 vssd1 vccd1 vccd1 _17380_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_81_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16933_ _18764_/Q _16965_/A2 _16965_/B1 input229/X _16965_/C1 vssd1 vssd1 vccd1 vccd1
+ _16933_/X sky130_fd_sc_hd__a221o_4
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12056_ _09494_/A _12086_/A2 _12055_/X _14340_/A vssd1 vssd1 vccd1 vccd1 _17805_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_238_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1831 _17326_/A vssd1 vssd1 vccd1 vccd1 _17338_/A sky130_fd_sc_hd__buf_4
Xfanout1842 _12428_/C1 vssd1 vssd1 vccd1 vccd1 _14181_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_237_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1853 _16960_/A vssd1 vssd1 vccd1 vccd1 _16904_/A sky130_fd_sc_hd__buf_2
XFILLER_238_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11007_ _19053_/Q _19021_/Q _11395_/C vssd1 vssd1 vccd1 vccd1 _11007_/X sky130_fd_sc_hd__mux2_1
Xfanout1864 _16964_/A vssd1 vssd1 vccd1 vccd1 _16972_/A sky130_fd_sc_hd__buf_4
XFILLER_38_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19652_ _19652_/A vssd1 vssd1 vccd1 vccd1 _19652_/X sky130_fd_sc_hd__buf_2
Xfanout1875 _17261_/A vssd1 vssd1 vccd1 vccd1 _17231_/A sky130_fd_sc_hd__buf_6
X_16864_ _18747_/Q _12276_/A _16877_/B1 input242/X _08828_/A vssd1 vssd1 vccd1 vccd1
+ _16864_/X sky130_fd_sc_hd__a221o_1
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1886 fanout1905/X vssd1 vssd1 vccd1 vccd1 _17725_/C1 sky130_fd_sc_hd__buf_6
XFILLER_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1897 _16110_/B1 vssd1 vssd1 vccd1 vccd1 _16737_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_237_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18603_ _19595_/CLK _18603_/D vssd1 vssd1 vccd1 vccd1 _18603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15815_ _18607_/Q _17705_/A0 _15832_/S vssd1 vssd1 vccd1 vccd1 _18607_/D sky130_fd_sc_hd__mux2_1
XFILLER_237_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19583_ _19615_/CLK _19583_/D vssd1 vssd1 vccd1 vccd1 _19583_/Q sky130_fd_sc_hd__dfxtp_1
X_16795_ _16795_/A _16795_/B _16799_/C vssd1 vssd1 vccd1 vccd1 _19286_/D sky130_fd_sc_hd__nor3_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15746_ _18591_/Q _18590_/Q _15746_/C vssd1 vssd1 vccd1 vccd1 _15772_/B sky130_fd_sc_hd__and3_1
X_18534_ _19620_/CLK _18534_/D vssd1 vssd1 vccd1 vccd1 _18534_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12958_ _13224_/B _14141_/D _12956_/X _13227_/C1 vssd1 vssd1 vccd1 vccd1 _12958_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_240_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11909_ _11909_/A _11909_/B vssd1 vssd1 vccd1 vccd1 _11909_/X sky130_fd_sc_hd__and2_1
XFILLER_206_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15677_ _18588_/Q _15704_/C vssd1 vssd1 vccd1 vccd1 _15677_/Y sky130_fd_sc_hd__nand2_1
X_18465_ _19644_/CLK _18465_/D vssd1 vssd1 vccd1 vccd1 _18465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12889_ _12883_/Y _12888_/Y _13263_/A vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__mux2_1
XANTENNA_270 input230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_281 input244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14628_ _16488_/A0 _18435_/Q _14628_/S vssd1 vssd1 vccd1 vccd1 _18435_/D sky130_fd_sc_hd__mux2_1
XANTENNA_292 _11922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17416_ _18567_/Q _17461_/A2 _17546_/A2 vssd1 vssd1 vccd1 vccd1 _17416_/X sky130_fd_sc_hd__o21a_1
XFILLER_159_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18396_ _19399_/CLK _18396_/D vssd1 vssd1 vccd1 vccd1 _18396_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_187_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17347_ _19471_/Q _17589_/A _17361_/S vssd1 vssd1 vccd1 vccd1 _17348_/B sky130_fd_sc_hd__mux2_1
X_14559_ _18388_/Q _14559_/A2 _14559_/B1 input16/X vssd1 vssd1 vccd1 vccd1 _14560_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17278_ _18120_/Q _15782_/A1 _17488_/A _17289_/B vssd1 vssd1 vccd1 vccd1 _17278_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_228_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16229_ _17693_/A0 _18844_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _18844_/D sky130_fd_sc_hd__mux2_1
X_19017_ _19216_/CLK _19017_/D vssd1 vssd1 vccd1 vccd1 _19017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08982_ _08980_/X _08981_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _08982_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09603_ _10366_/A1 _18209_/Q _09720_/S _18944_/Q _10371_/S vssd1 vssd1 vccd1 vccd1
+ _09603_/X sky130_fd_sc_hd__o221a_1
XFILLER_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09534_ _09532_/X _09533_/X _09534_/S vssd1 vssd1 vccd1 vccd1 _09535_/B sky130_fd_sc_hd__mux2_1
XFILLER_225_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09465_ _10263_/A1 _18140_/Q _18786_/Q _09464_/S vssd1 vssd1 vccd1 vccd1 _09465_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09396_ _11046_/S1 _09386_/X _09395_/X _11438_/B1 vssd1 vssd1 vccd1 vccd1 _09396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_212_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_173_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19542_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_102_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18715_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10240_ _18467_/Q _18368_/Q _10253_/C vssd1 vssd1 vccd1 vccd1 _10240_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ _11017_/A1 _19224_/Q _19192_/Q _10176_/S _11397_/A1 vssd1 vssd1 vccd1 vccd1
+ _10171_/X sky130_fd_sc_hd__a221o_1
XFILLER_65_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput480 _18109_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[8] sky130_fd_sc_hd__buf_4
XFILLER_267_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1105 _12589_/X vssd1 vssd1 vccd1 vccd1 _13563_/B1 sky130_fd_sc_hd__buf_4
Xfanout1116 _13941_/B vssd1 vssd1 vccd1 vccd1 _13818_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1127 _15140_/B vssd1 vssd1 vccd1 vccd1 _15411_/B sky130_fd_sc_hd__buf_4
Xfanout1138 _16500_/A0 vssd1 vssd1 vccd1 vccd1 _17666_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1149 _09103_/Y vssd1 vssd1 vccd1 vccd1 _11024_/A1 sky130_fd_sc_hd__buf_8
XFILLER_87_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13930_ _13930_/A1 _13917_/Y _13930_/B1 vssd1 vssd1 vccd1 vccd1 _13931_/C sky130_fd_sc_hd__o21a_1
XFILLER_275_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13861_ _13861_/A _14150_/B vssd1 vssd1 vccd1 vccd1 _13861_/Y sky130_fd_sc_hd__nand2_1
XFILLER_207_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15600_ _15580_/A _15580_/B _15577_/X _15576_/X vssd1 vssd1 vccd1 vccd1 _15602_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_170_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12812_ _12703_/X _12712_/X _12813_/S vssd1 vssd1 vccd1 vccd1 _12812_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16580_ _16580_/A0 _19184_/Q _16585_/S vssd1 vssd1 vccd1 vccd1 _19184_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13792_ _13622_/A _13807_/B _13323_/X _13791_/X vssd1 vssd1 vccd1 vccd1 _13792_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_62_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15531_ _15531_/A _15531_/B vssd1 vssd1 vccd1 vccd1 _15554_/B sky130_fd_sc_hd__xnor2_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12743_/A _13961_/A vssd1 vssd1 vccd1 vccd1 _12746_/B sky130_fd_sc_hd__nor2_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _19632_/CLK _18250_/D vssd1 vssd1 vccd1 vccd1 _18250_/Q sky130_fd_sc_hd__dfxtp_1
X_15462_ _15557_/A _15558_/A vssd1 vssd1 vccd1 vccd1 _15464_/A sky130_fd_sc_hd__and2_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12673_/X _12672_/Y _12818_/S vssd1 vssd1 vccd1 vccd1 _12674_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17210_/A _17201_/B vssd1 vssd1 vccd1 vccd1 _19418_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14413_ _16455_/A1 _18264_/Q _14415_/S vssd1 vssd1 vccd1 vccd1 _18264_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18181_ _19634_/CLK _18181_/D vssd1 vssd1 vccd1 vccd1 _18181_/Q sky130_fd_sc_hd__dfxtp_1
X_11625_ _14268_/A _13941_/A _13904_/A vssd1 vssd1 vccd1 vccd1 _13962_/A sky130_fd_sc_hd__mux2_8
XFILLER_168_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15393_ _15223_/A _15390_/Y _15392_/Y _15416_/A vssd1 vssd1 vccd1 vccd1 _15393_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_11_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17132_ _19395_/Q _17120_/Y _17131_/X vssd1 vssd1 vccd1 vccd1 _19395_/D sky130_fd_sc_hd__o21ba_1
X_14344_ _15039_/A _14345_/B _14344_/C vssd1 vssd1 vccd1 vccd1 _18199_/D sky130_fd_sc_hd__and3_4
XFILLER_200_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11556_ _11556_/A _11556_/B _11556_/C vssd1 vssd1 vccd1 vccd1 _11556_/X sky130_fd_sc_hd__or3_1
XFILLER_155_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17063_ _19365_/Q _17113_/B vssd1 vssd1 vccd1 vccd1 _17063_/X sky130_fd_sc_hd__or2_1
X_10507_ _18619_/Q _18190_/Q _10511_/S vssd1 vssd1 vccd1 vccd1 _10507_/X sky130_fd_sc_hd__mux2_1
X_14275_ _17693_/A0 _18134_/Q _14277_/S vssd1 vssd1 vccd1 vccd1 _18134_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11487_ _10239_/A _11486_/X _11452_/Y _11790_/B vssd1 vssd1 vccd1 vccd1 _11819_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_171_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16014_ _18722_/Q _16016_/A2 _16147_/A2 _18771_/Q _16018_/C1 vssd1 vssd1 vccd1 vccd1
+ _16014_/X sky130_fd_sc_hd__a221o_1
X_13226_ _13226_/A _13226_/B vssd1 vssd1 vccd1 vccd1 _13226_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ _11596_/A1 _18159_/Q _18805_/Q _10815_/B vssd1 vssd1 vccd1 vccd1 _10438_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13157_ _13896_/B2 _13153_/X _13156_/Y _12732_/S _13155_/Y vssd1 vssd1 vccd1 vccd1
+ _13157_/X sky130_fd_sc_hd__o221a_4
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10369_ _18466_/Q _18367_/Q _10370_/S vssd1 vssd1 vccd1 vccd1 _10369_/X sky130_fd_sc_hd__mux2_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _17829_/Q _12104_/B _12107_/Y vssd1 vssd1 vccd1 vccd1 _17829_/D sky130_fd_sc_hd__o21a_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _17982_/CLK _17965_/D vssd1 vssd1 vccd1 vccd1 _17965_/Q sky130_fd_sc_hd__dfxtp_1
X_13088_ _13086_/X _13087_/X _13135_/S vssd1 vssd1 vccd1 vccd1 _13088_/X sky130_fd_sc_hd__mux2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16916_ _16928_/A _16916_/B vssd1 vssd1 vccd1 vccd1 _19313_/D sky130_fd_sc_hd__and2_1
Xfanout1650 _09873_/A1 vssd1 vssd1 vccd1 vccd1 _08901_/A sky130_fd_sc_hd__buf_8
X_12039_ _17797_/Q _12051_/B vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__or2_1
Xfanout1661 _09873_/A1 vssd1 vssd1 vccd1 vccd1 _11498_/A1 sky130_fd_sc_hd__buf_6
Xfanout1672 _10746_/S vssd1 vssd1 vccd1 vccd1 _10301_/S sky130_fd_sc_hd__buf_12
X_17896_ _18817_/CLK _17896_/D vssd1 vssd1 vccd1 vccd1 _17896_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1683 _09854_/A vssd1 vssd1 vccd1 vccd1 _11157_/A1 sky130_fd_sc_hd__buf_6
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1694 _11404_/A1 vssd1 vssd1 vccd1 vccd1 _10334_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_238_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19635_ _19635_/CLK _19635_/D vssd1 vssd1 vccd1 vccd1 _19635_/Q sky130_fd_sc_hd__dfxtp_1
X_16847_ _19296_/Q _16967_/S _16846_/Y _16968_/A vssd1 vssd1 vccd1 vccd1 _19296_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19566_ _19612_/CLK _19566_/D vssd1 vssd1 vccd1 vccd1 _19566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16778_ _19280_/Q _16778_/B vssd1 vssd1 vccd1 vccd1 _16783_/C sky130_fd_sc_hd__and2_2
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18517_ _18517_/CLK _18517_/D vssd1 vssd1 vccd1 vccd1 _18517_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_207_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15729_ _18590_/Q _15746_/C vssd1 vssd1 vccd1 vccd1 _15729_/X sky130_fd_sc_hd__and2_1
XFILLER_234_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_0_wb_clk_i _19652_/A vssd1 vssd1 vccd1 vccd1 _19632_/CLK sky130_fd_sc_hd__clkbuf_16
X_19497_ _19533_/CLK _19497_/D vssd1 vssd1 vccd1 vccd1 _19497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09250_ _18852_/Q _18884_/Q _09269_/S vssd1 vssd1 vccd1 vccd1 _09250_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18448_ _19627_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09181_ _19077_/Q _18981_/Q _09181_/S vssd1 vssd1 vccd1 vccd1 _09181_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18379_ _19465_/CLK _18379_/D vssd1 vssd1 vccd1 vccd1 _18379_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_119_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08965_ _11497_/A1 _19206_/Q _19174_/Q _09952_/S vssd1 vssd1 vccd1 vccd1 _08965_/X
+ sky130_fd_sc_hd__a22o_1
Xinput208 localMemory_wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__clkbuf_2
Xinput219 localMemory_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input219/X sky130_fd_sc_hd__buf_8
XFILLER_69_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08896_ _08896_/A _09285_/C vssd1 vssd1 vccd1 vccd1 _08896_/Y sky130_fd_sc_hd__nand2_2
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09517_ _19073_/Q _18977_/Q _09883_/B vssd1 vssd1 vccd1 vccd1 _09517_/X sky130_fd_sc_hd__mux2_1
XFILLER_225_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _10266_/S1 _09447_/X _09446_/X _09463_/S vssd1 vssd1 vccd1 vccd1 _09448_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09379_ _18447_/Q _18348_/Q _10141_/S vssd1 vssd1 vccd1 vccd1 _09379_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11410_ _10239_/A _11409_/Y _11376_/Y _11790_/B vssd1 vssd1 vccd1 vccd1 _11823_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_137_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ _18390_/Q _12429_/B1 _09236_/Y _08858_/A vssd1 vssd1 vccd1 vccd1 _12391_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_137_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11341_ _11339_/X _11340_/X _11361_/S vssd1 vssd1 vccd1 vccd1 _11341_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ _17677_/A0 _18002_/Q _14072_/S vssd1 vssd1 vccd1 vccd1 _18002_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11272_ _11282_/A _11271_/X _11286_/B1 vssd1 vssd1 vccd1 vccd1 _11272_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13011_ _19237_/Q _13495_/A2 _13495_/B1 _19269_/Q vssd1 vssd1 vccd1 vccd1 _13011_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10223_ _18468_/Q _18369_/Q _10224_/S vssd1 vssd1 vccd1 vccd1 _10223_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_70_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19612_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10154_ _10147_/X _10153_/X _10137_/X vssd1 vssd1 vccd1 vccd1 _10154_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_160_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14962_ _17817_/Q _14982_/B vssd1 vssd1 vccd1 vccd1 _14962_/X sky130_fd_sc_hd__or2_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17750_ _18650_/Q vssd1 vssd1 vccd1 vccd1 _18650_/D sky130_fd_sc_hd__clkbuf_2
X_10085_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10309_/B sky130_fd_sc_hd__nand2_2
XFILLER_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16701_ _19253_/Q _16704_/C vssd1 vssd1 vccd1 vccd1 _16701_/Y sky130_fd_sc_hd__nand2_1
XFILLER_248_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13913_ _13913_/A _13913_/B vssd1 vssd1 vccd1 vccd1 _13913_/X sky130_fd_sc_hd__or2_1
X_17681_ _17681_/A0 _19608_/Q _17681_/S vssd1 vssd1 vccd1 vccd1 _19608_/D sky130_fd_sc_hd__mux2_1
X_14893_ _18121_/Q _14892_/X _14893_/S vssd1 vssd1 vccd1 vccd1 _14893_/X sky130_fd_sc_hd__mux2_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19420_ _19485_/CLK _19420_/D vssd1 vssd1 vccd1 vccd1 _19420_/Q sky130_fd_sc_hd__dfxtp_1
X_16632_ _17724_/A _19232_/Q _19233_/Q vssd1 vssd1 vccd1 vccd1 _16634_/B sky130_fd_sc_hd__a21oi_1
X_13844_ _17851_/Q _13844_/A2 _13844_/B1 _17883_/Q vssd1 vssd1 vccd1 vccd1 _13844_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19351_ _19481_/CLK _19351_/D vssd1 vssd1 vccd1 vccd1 _19351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16563_ _17696_/A0 _19167_/Q _16586_/S vssd1 vssd1 vccd1 vccd1 _19167_/D sky130_fd_sc_hd__mux2_1
X_13775_ _13775_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13775_/X sky130_fd_sc_hd__or2_1
XFILLER_222_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ _17970_/Q _11447_/A2 _11371_/B1 vssd1 vssd1 vccd1 vccd1 _10988_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18302_ _19450_/CLK _18302_/D vssd1 vssd1 vccd1 vccd1 _18302_/Q sky130_fd_sc_hd__dfxtp_1
X_12726_ _12726_/A vssd1 vssd1 vccd1 vccd1 _12726_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15514_ _15561_/C _15514_/B vssd1 vssd1 vccd1 vccd1 _15514_/Y sky130_fd_sc_hd__nor2_1
X_19282_ _19285_/CLK _19282_/D vssd1 vssd1 vccd1 vccd1 _19282_/Q sky130_fd_sc_hd__dfxtp_1
X_16494_ _17660_/A0 _19100_/Q _16521_/S vssd1 vssd1 vccd1 vccd1 _19100_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18233_ _19613_/CLK _18233_/D vssd1 vssd1 vccd1 vccd1 _18233_/Q sky130_fd_sc_hd__dfxtp_1
X_15445_ _15445_/A _15445_/B vssd1 vssd1 vccd1 vccd1 _15445_/Y sky130_fd_sc_hd__xnor2_1
X_12657_ _10233_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _12657_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_157_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11608_ _08874_/D _11607_/X _11602_/X _11608_/C1 vssd1 vssd1 vccd1 vccd1 _11608_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_198_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18164_ _19607_/CLK _18164_/D vssd1 vssd1 vccd1 vccd1 _18164_/Q sky130_fd_sc_hd__dfxtp_1
X_15376_ _15376_/A _15376_/B vssd1 vssd1 vccd1 vccd1 _15376_/X sky130_fd_sc_hd__xor2_1
X_12588_ _12754_/B _12455_/A _12587_/B vssd1 vssd1 vccd1 vccd1 _12588_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_11_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17115_ _19391_/Q _17115_/B vssd1 vssd1 vccd1 vccd1 _17115_/X sky130_fd_sc_hd__or2_1
X_14327_ _18184_/Q _17678_/A0 _14339_/S vssd1 vssd1 vccd1 vccd1 _18184_/D sky130_fd_sc_hd__mux2_1
X_18095_ _18761_/CLK _18095_/D vssd1 vssd1 vccd1 vccd1 _18095_/Q sky130_fd_sc_hd__dfxtp_1
X_11539_ _12638_/A _11669_/B _10754_/A vssd1 vssd1 vccd1 vccd1 _11667_/A sky130_fd_sc_hd__a21o_2
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17046_ _17214_/B _17046_/A2 _17045_/X _17354_/A vssd1 vssd1 vccd1 vccd1 _19359_/D
+ sky130_fd_sc_hd__o211a_1
X_14258_ _18127_/Q _14260_/B vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__or2_1
XFILLER_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ _19499_/Q _13781_/A2 _13781_/B1 _13208_/X vssd1 vssd1 vccd1 vccd1 _13209_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14189_ _16972_/A _14189_/B vssd1 vssd1 vccd1 vccd1 _18092_/D sky130_fd_sc_hd__and2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout909 _16421_/S vssd1 vssd1 vccd1 vccd1 _16424_/S sky130_fd_sc_hd__buf_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _19157_/CLK _18997_/D vssd1 vssd1 vccd1 vccd1 _18997_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17948_ _18749_/CLK _17948_/D vssd1 vssd1 vccd1 vccd1 _17948_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1480 fanout1485/X vssd1 vssd1 vccd1 vccd1 _09801_/S sky130_fd_sc_hd__buf_4
Xfanout1491 _10721_/S vssd1 vssd1 vccd1 vccd1 _10362_/S sky130_fd_sc_hd__buf_6
XFILLER_66_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17879_ _19320_/CLK _17879_/D vssd1 vssd1 vccd1 vccd1 _17879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19618_ _19618_/CLK _19618_/D vssd1 vssd1 vccd1 vccd1 _19618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19549_ _19553_/CLK _19549_/D vssd1 vssd1 vccd1 vccd1 _19549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09302_ _18025_/Q _17993_/Q _09302_/S vssd1 vssd1 vccd1 vccd1 _09302_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09233_ _18398_/Q _09656_/B1 _09232_/Y _09992_/A vssd1 vssd1 vccd1 vccd1 _09902_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_142_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09164_ _18542_/Q _18417_/Q _09179_/B vssd1 vssd1 vccd1 vccd1 _09164_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09095_ _09095_/A _12023_/A vssd1 vssd1 vccd1 vccd1 _09095_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_2__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_266_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ _11157_/A1 _17758_/Q _11226_/S _18307_/Q _11567_/S vssd1 vssd1 vccd1 vccd1
+ _09997_/X sky130_fd_sc_hd__o221a_1
XFILLER_135_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _08948_/A _08948_/B vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__nand2_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ _12460_/A _12320_/A _10471_/S _12320_/B vssd1 vssd1 vccd1 vccd1 _08880_/D
+ sky130_fd_sc_hd__or4_2
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ _10085_/A _09037_/X _11143_/A1 vssd1 vssd1 vccd1 vccd1 _10912_/A sky130_fd_sc_hd__a21oi_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _11899_/A _11890_/B _11890_/C vssd1 vssd1 vccd1 vccd1 _11890_/X sky130_fd_sc_hd__and3_4
XFILLER_260_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _11562_/S _10840_/X _10839_/X _10841_/C1 vssd1 vssd1 vccd1 vccd1 _10841_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_260_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13560_ _13682_/B2 _13549_/X _13551_/Y _13559_/Y vssd1 vssd1 vccd1 vccd1 _14012_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_13_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10772_ _11327_/S _18800_/Q _10856_/C vssd1 vssd1 vccd1 vccd1 _10772_/X sky130_fd_sc_hd__and3_1
XFILLER_213_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _12553_/A _12553_/B _12553_/C _12553_/D vssd1 vssd1 vccd1 vccd1 _12512_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_201_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13491_ _13622_/A _13512_/B vssd1 vssd1 vccd1 vccd1 _13491_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15230_ _15228_/Y _15230_/B vssd1 vssd1 vccd1 vccd1 _15233_/A sky130_fd_sc_hd__and2b_1
XFILLER_185_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _12442_/A _12442_/B _12442_/C _12442_/D vssd1 vssd1 vccd1 vccd1 _12443_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15161_ _18565_/Q _18564_/Q vssd1 vssd1 vccd1 vccd1 _15161_/Y sky130_fd_sc_hd__xnor2_1
X_12373_ _12427_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _12373_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14112_ _16529_/A0 _18051_/Q _14140_/S vssd1 vssd1 vccd1 vccd1 _18051_/D sky130_fd_sc_hd__mux2_1
X_11324_ _11322_/X _11323_/X _11577_/S vssd1 vssd1 vccd1 vccd1 _11324_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15092_ _19379_/Q _15092_/B _15092_/C vssd1 vssd1 vccd1 vccd1 _15092_/X sky130_fd_sc_hd__and3_1
XFILLER_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18920_ _19631_/CLK _18920_/D vssd1 vssd1 vccd1 vccd1 _18920_/Q sky130_fd_sc_hd__dfxtp_1
X_14043_ _16593_/A0 _17985_/Q _14070_/S vssd1 vssd1 vccd1 vccd1 _17985_/D sky130_fd_sc_hd__mux2_1
X_11255_ _09086_/A _11252_/X _11245_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _11255_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_268_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10206_ _19096_/Q _19000_/Q _10206_/S vssd1 vssd1 vccd1 vccd1 _10206_/X sky130_fd_sc_hd__mux2_1
X_18851_ _19626_/CLK _18851_/D vssd1 vssd1 vccd1 vccd1 _18851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11186_ _11184_/X _11185_/X _11198_/S vssd1 vssd1 vccd1 vccd1 _11186_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17802_ _19650_/CLK _17802_/D vssd1 vssd1 vccd1 vccd1 _17802_/Q sky130_fd_sc_hd__dfxtp_4
X_10137_ _11053_/A _10131_/X _10134_/X _10136_/X _11417_/B1 vssd1 vssd1 vccd1 vccd1
+ _10137_/X sky130_fd_sc_hd__a311o_2
XFILLER_39_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18782_ _19589_/CLK _18782_/D vssd1 vssd1 vccd1 vccd1 _18782_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15994_ _18712_/Q _16002_/A2 _16002_/B1 _18761_/Q _16002_/C1 vssd1 vssd1 vccd1 vccd1
+ _15994_/X sky130_fd_sc_hd__a221o_1
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17733_ _18633_/Q vssd1 vssd1 vccd1 vccd1 _18633_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_36_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10068_ _11731_/B _10068_/B vssd1 vssd1 vccd1 vccd1 _11735_/A sky130_fd_sc_hd__nand2_2
X_14945_ _18126_/Q _14893_/S _14934_/X _14944_/X vssd1 vssd1 vccd1 vccd1 _14945_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17664_ _17664_/A0 _19591_/Q _17687_/S vssd1 vssd1 vccd1 vccd1 _19591_/D sky130_fd_sc_hd__mux2_1
XFILLER_235_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14876_ input52/X input88/X _14947_/S vssd1 vssd1 vccd1 vccd1 _14877_/A sky130_fd_sc_hd__mux2_2
X_19403_ _19466_/CLK _19403_/D vssd1 vssd1 vccd1 vccd1 _19403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16615_ _16615_/A0 _19218_/Q _16618_/S vssd1 vssd1 vccd1 vccd1 _19218_/D sky130_fd_sc_hd__mux2_1
X_13827_ _19355_/Q _13883_/A2 _13883_/B1 _19483_/Q _13883_/C1 vssd1 vssd1 vccd1 vccd1
+ _13827_/X sky130_fd_sc_hd__a221o_1
X_17595_ _19377_/Q _15086_/B input178/X _17592_/X _17623_/B1 vssd1 vssd1 vccd1 vccd1
+ _17595_/X sky130_fd_sc_hd__a41o_1
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19334_ _19534_/CLK _19334_/D vssd1 vssd1 vccd1 vccd1 _19334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13758_ _13758_/A _13758_/B vssd1 vssd1 vccd1 vccd1 _13758_/Y sky130_fd_sc_hd__nand2_1
X_16546_ _17679_/A0 _19151_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _19151_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12709_ _12707_/X _12708_/X _12813_/S vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__mux2_1
X_19265_ _19268_/CLK _19265_/D vssd1 vssd1 vccd1 vccd1 _19265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13689_ _19383_/Q _13884_/A2 _13687_/X _13688_/X _13884_/C1 vssd1 vssd1 vccd1 vccd1
+ _13689_/X sky130_fd_sc_hd__o221a_4
X_16477_ _16543_/A0 _19084_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _19084_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18216_ _19612_/CLK _18216_/D vssd1 vssd1 vccd1 vccd1 _18216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15428_ _18116_/Q _15133_/Y _15427_/X _15429_/A2 vssd1 vssd1 vccd1 vccd1 _15432_/A
+ sky130_fd_sc_hd__a22o_2
X_19196_ _19196_/CLK _19196_/D vssd1 vssd1 vccd1 vccd1 _19196_/Q sky130_fd_sc_hd__dfxtp_1
X_18147_ _19216_/CLK _18147_/D vssd1 vssd1 vccd1 vccd1 _18147_/Q sky130_fd_sc_hd__dfxtp_1
X_15359_ _18113_/Q _15132_/X _15358_/X _15429_/A2 vssd1 vssd1 vccd1 vccd1 _15361_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_129_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18078_ _19628_/CLK _18078_/D vssd1 vssd1 vccd1 vccd1 _18078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09920_ _10262_/A1 _19132_/Q _11472_/C _19100_/Q _09935_/A vssd1 vssd1 vccd1 vccd1
+ _09920_/X sky130_fd_sc_hd__o221a_1
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17029_ _19351_/Q _17041_/B vssd1 vssd1 vccd1 vccd1 _17029_/X sky130_fd_sc_hd__or2_1
Xfanout706 _12543_/X vssd1 vssd1 vccd1 vccd1 _13821_/B sky130_fd_sc_hd__clkbuf_4
Xfanout717 _13952_/A2 vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__buf_8
XFILLER_59_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09851_ _18018_/Q _17986_/Q _10001_/S vssd1 vssd1 vccd1 vccd1 _09851_/X sky130_fd_sc_hd__mux2_1
Xfanout728 _16538_/A0 vssd1 vssd1 vccd1 vccd1 _17704_/A0 sky130_fd_sc_hd__buf_4
XFILLER_140_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout739 _11299_/X vssd1 vssd1 vccd1 vccd1 _16507_/A0 sky130_fd_sc_hd__buf_2
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09782_ _19038_/Q _19006_/Q _09797_/S vssd1 vssd1 vccd1 vccd1 _09782_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09216_ _19109_/Q _19141_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _09216_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09147_ _09908_/A1 _09232_/A _09146_/X _09908_/B1 _18399_/Q vssd1 vssd1 vccd1 vccd1
+ _09819_/C sky130_fd_sc_hd__o32a_1
XFILLER_136_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ _17894_/Q _17893_/Q _17892_/Q _09062_/B vssd1 vssd1 vccd1 vccd1 _09080_/C
+ sky130_fd_sc_hd__o31a_2
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11040_ _11498_/A1 _19213_/Q _19181_/Q _09966_/S vssd1 vssd1 vccd1 vccd1 _11040_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _13046_/A1 _12989_/Y _12990_/X vssd1 vssd1 vccd1 vccd1 _12992_/A sky130_fd_sc_hd__o21ai_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14730_ _14727_/Y _14729_/Y _14950_/B1 vssd1 vssd1 vccd1 vccd1 _14730_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_55_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11942_ _11944_/A1 _11868_/B _11959_/A2 input229/X vssd1 vssd1 vccd1 vccd1 _11942_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14661_ _17720_/A0 _18467_/Q _14663_/S vssd1 vssd1 vccd1 vccd1 _18467_/D sky130_fd_sc_hd__mux2_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11873_ _10564_/B _11864_/B _11926_/A1 vssd1 vssd1 vccd1 vccd1 _11878_/B sky130_fd_sc_hd__o21ai_2
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16400_ _17665_/A0 _19009_/Q _16421_/S vssd1 vssd1 vccd1 vccd1 _19009_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13612_ _10027_/A _13971_/A2 _13610_/Y _13611_/X _13579_/A vssd1 vssd1 vccd1 vccd1
+ _13612_/X sky130_fd_sc_hd__a221o_4
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10824_ _10822_/X _10823_/X _11601_/A vssd1 vssd1 vccd1 vccd1 _10824_/X sky130_fd_sc_hd__mux2_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14592_ _14592_/A _14592_/B vssd1 vssd1 vccd1 vccd1 _18404_/D sky130_fd_sc_hd__or2_1
X_17380_ _17380_/A _17380_/B vssd1 vssd1 vccd1 vccd1 _19487_/D sky130_fd_sc_hd__and2_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16331_ _18943_/Q _17663_/A0 _16355_/S vssd1 vssd1 vccd1 vccd1 _18943_/D sky130_fd_sc_hd__mux2_1
X_13543_ _15452_/A _13539_/X _13542_/X _13869_/B2 vssd1 vssd1 vccd1 vccd1 _13544_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10755_ _12638_/A vssd1 vssd1 vccd1 vccd1 _13665_/A sky130_fd_sc_hd__clkinv_2
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16262_ _17693_/A0 _18876_/Q _16288_/S vssd1 vssd1 vccd1 vccd1 _18876_/D sky130_fd_sc_hd__mux2_1
X_19050_ _19640_/CLK _19050_/D vssd1 vssd1 vccd1 vccd1 _19050_/Q sky130_fd_sc_hd__dfxtp_1
X_13474_ _13899_/A _13472_/X _13473_/Y _13970_/B2 vssd1 vssd1 vccd1 vccd1 _13475_/B
+ sky130_fd_sc_hd__a22o_1
X_10686_ _11250_/A1 _19217_/Q _19185_/Q _10687_/S _11480_/C1 vssd1 vssd1 vccd1 vccd1
+ _10686_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18001_ _19148_/CLK _18001_/D vssd1 vssd1 vccd1 vccd1 _18001_/Q sky130_fd_sc_hd__dfxtp_1
X_15213_ _17914_/Q _15369_/A vssd1 vssd1 vccd1 vccd1 _15219_/A sky130_fd_sc_hd__nand2_2
X_12425_ _17916_/Q _12421_/A _12424_/Y _12428_/C1 vssd1 vssd1 vccd1 vccd1 _17916_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16193_ _16292_/A0 _18810_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _18810_/D sky130_fd_sc_hd__mux2_1
XFILLER_275_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15144_ _19458_/Q _19392_/Q _15400_/S vssd1 vssd1 vccd1 vccd1 _15145_/C sky130_fd_sc_hd__and3_1
X_12356_ _17893_/Q _12379_/A _12355_/Y _13981_/C1 vssd1 vssd1 vccd1 vccd1 _17893_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput309 _11757_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[13] sky130_fd_sc_hd__buf_4
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11307_ _18546_/Q _11309_/S vssd1 vssd1 vccd1 vccd1 _11307_/X sky130_fd_sc_hd__or2_1
X_15075_ _18559_/Q _17686_/A0 _15078_/S vssd1 vssd1 vccd1 vccd1 _18559_/D sky130_fd_sc_hd__mux2_1
XFILLER_236_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12287_ _18088_/Q _12305_/A2 _12305_/B1 _18511_/Q vssd1 vssd1 vccd1 vccd1 _12486_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18903_ _19614_/CLK _18903_/D vssd1 vssd1 vccd1 vccd1 _18903_/Q sky130_fd_sc_hd__dfxtp_1
X_14026_ _14028_/A _14026_/B vssd1 vssd1 vccd1 vccd1 _14026_/Y sky130_fd_sc_hd__nand2_1
X_11238_ _18454_/Q _18355_/Q _11247_/S vssd1 vssd1 vccd1 vccd1 _11238_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18834_ _19644_/CLK _18834_/D vssd1 vssd1 vccd1 vccd1 _18834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11169_ _11172_/A1 _18610_/Q _18181_/Q _11160_/S vssd1 vssd1 vccd1 vccd1 _11169_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18765_ _19076_/CLK _18765_/D vssd1 vssd1 vccd1 vccd1 _18765_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15977_ _18704_/Q _15977_/A2 _15976_/X _16972_/A vssd1 vssd1 vccd1 vccd1 _18704_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17716_ _17716_/A0 _19642_/Q _17718_/S vssd1 vssd1 vccd1 vccd1 _19642_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14928_ _14979_/A1 _18271_/Q _14927_/Y _14928_/B1 vssd1 vssd1 vccd1 vccd1 _14928_/X
+ sky130_fd_sc_hd__a31o_1
X_18696_ _19304_/CLK _18696_/D vssd1 vssd1 vccd1 vccd1 _18696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17647_ _17680_/A0 _19575_/Q _17657_/S vssd1 vssd1 vccd1 vccd1 _19575_/D sky130_fd_sc_hd__mux2_1
XFILLER_224_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14859_ _14855_/Y _14858_/X _14879_/B1 vssd1 vssd1 vccd1 vccd1 _14859_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17578_ _19531_/Q _17622_/A2 _17603_/B1 _17577_/X vssd1 vssd1 vccd1 vccd1 _19531_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19317_ _19502_/CLK _19317_/D vssd1 vssd1 vccd1 vccd1 _19317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16529_ _16529_/A0 _19134_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _19134_/D sky130_fd_sc_hd__mux2_1
X_19248_ _19268_/CLK _19248_/D vssd1 vssd1 vccd1 vccd1 _19248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09001_ _18268_/Q _18198_/Q vssd1 vssd1 vccd1 vccd1 _09652_/A sky130_fd_sc_hd__nand2_8
X_19179_ _19211_/CLK _19179_/D vssd1 vssd1 vccd1 vccd1 _19179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09903_ _11687_/A _09903_/B _09903_/C _09903_/D vssd1 vssd1 vccd1 vccd1 _09903_/X
+ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_198_wb_clk_i _19652_/A vssd1 vssd1 vccd1 vccd1 _19575_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout503 _11953_/B2 vssd1 vssd1 vccd1 vccd1 _11959_/B2 sky130_fd_sc_hd__buf_6
Xfanout514 _17289_/B vssd1 vssd1 vccd1 vccd1 _17307_/B sky130_fd_sc_hd__buf_4
XFILLER_98_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout525 _11899_/A vssd1 vssd1 vccd1 vccd1 _11818_/B sky130_fd_sc_hd__buf_4
Xfanout536 _17119_/X vssd1 vssd1 vccd1 vccd1 fanout536/X sky130_fd_sc_hd__buf_6
XFILLER_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_127_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19319_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout547 _15476_/A1 vssd1 vssd1 vccd1 vccd1 _17389_/B1 sky130_fd_sc_hd__buf_6
X_09834_ _09086_/A _09827_/X _09829_/X _09831_/X _09833_/X vssd1 vssd1 vccd1 vccd1
+ _09834_/X sky130_fd_sc_hd__o32a_1
XFILLER_258_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout558 _15764_/A vssd1 vssd1 vccd1 vccd1 _15787_/A sky130_fd_sc_hd__buf_6
XFILLER_247_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout569 _15113_/Y vssd1 vssd1 vccd1 vccd1 _15623_/A sky130_fd_sc_hd__buf_12
XFILLER_247_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09765_ _18629_/Q _18051_/Q _19070_/Q _18974_/Q _11226_/S _11569_/S1 vssd1 vssd1
+ vccd1 vccd1 _09765_/X sky130_fd_sc_hd__mux4_1
XFILLER_274_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09696_ _15120_/A _11793_/B _09695_/Y _10027_/B vssd1 vssd1 vccd1 vccd1 _09696_/X
+ sky130_fd_sc_hd__a211o_2
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10540_ _11583_/A _10539_/Y _10536_/Y _09086_/A vssd1 vssd1 vccd1 vccd1 _10540_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10471_ _10469_/X _10470_/X _10471_/S vssd1 vssd1 vccd1 vccd1 _10471_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12210_ _17868_/Q _12210_/B vssd1 vssd1 vccd1 vccd1 _12216_/C sky130_fd_sc_hd__and2_2
XFILLER_136_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13190_ _13349_/B _14143_/C _13260_/A vssd1 vssd1 vccd1 vccd1 _13190_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12141_ _17842_/Q _12144_/C _17330_/A vssd1 vssd1 vccd1 vccd1 _12141_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12072_ _09777_/A _12086_/A2 _12071_/X _17419_/C1 vssd1 vssd1 vccd1 vccd1 _17813_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15900_ _18675_/Q _15906_/A2 _15903_/B1 _15899_/X vssd1 vssd1 vccd1 vccd1 _15900_/X
+ sky130_fd_sc_hd__a211o_1
X_11023_ _11452_/A _16610_/A0 _11023_/B1 vssd1 vssd1 vccd1 vccd1 _11023_/X sky130_fd_sc_hd__o21a_1
XFILLER_173_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16880_ _16968_/A _16880_/B vssd1 vssd1 vccd1 vccd1 _19304_/D sky130_fd_sc_hd__and2_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15831_ _18623_/Q _16621_/A0 _15832_/S vssd1 vssd1 vccd1 vccd1 _18623_/D sky130_fd_sc_hd__mux2_1
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18550_ _19636_/CLK _18550_/D vssd1 vssd1 vccd1 vccd1 _18550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ input5/X _12552_/X _12967_/X _12973_/X _12538_/B vssd1 vssd1 vccd1 vccd1
+ _12974_/X sky130_fd_sc_hd__o221a_2
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _13935_/Y _15110_/X _10156_/Y _15502_/B vssd1 vssd1 vccd1 vccd1 _15762_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _18584_/Q _17544_/A _17516_/C1 vssd1 vssd1 vccd1 vccd1 _17501_/X sky130_fd_sc_hd__o21a_1
XFILLER_261_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _17792_/Q _14712_/X _14993_/S vssd1 vssd1 vccd1 vccd1 _14713_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18481_ _18517_/CLK _18481_/D vssd1 vssd1 vccd1 vccd1 _18481_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11925_ _11926_/A1 _11939_/A1 _11825_/B _11935_/B1 input242/X vssd1 vssd1 vccd1 vccd1
+ _11925_/X sky130_fd_sc_hd__a32o_4
XFILLER_46_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _19482_/Q _19416_/Q vssd1 vssd1 vccd1 vccd1 _15693_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_430 _11836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_441 _13996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_452 _14599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _18109_/Q _17437_/A2 _17430_/X _17431_/X vssd1 vssd1 vccd1 vccd1 _17432_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_261_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14644_ _16471_/A0 _18450_/Q _14663_/S vssd1 vssd1 vccd1 vccd1 _18450_/D sky130_fd_sc_hd__mux2_1
XFILLER_221_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_463 _18384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11856_ _11952_/A2 _11854_/X _11855_/X vssd1 vssd1 vccd1 vccd1 _11857_/B sky130_fd_sc_hd__a21oi_4
XFILLER_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_474 input222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_485 _11928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_496 _16589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ _11358_/A _10799_/X _10798_/X _11361_/S vssd1 vssd1 vccd1 vccd1 _10807_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17363_ _19479_/Q _17190_/B _17379_/S vssd1 vssd1 vccd1 vccd1 _17364_/B sky130_fd_sc_hd__mux2_1
X_14575_ _18396_/Q _14575_/A2 _14575_/B1 input25/X vssd1 vssd1 vccd1 vccd1 _14576_/B
+ sky130_fd_sc_hd__o22a_1
X_11787_ _11799_/A _11799_/B _11807_/B vssd1 vssd1 vccd1 vccd1 _11787_/X sky130_fd_sc_hd__and3_1
XFILLER_186_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19102_ _19134_/CLK _19102_/D vssd1 vssd1 vccd1 vccd1 _19102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16314_ _16314_/A0 _18927_/Q _16320_/S vssd1 vssd1 vccd1 vccd1 _18927_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13526_ _19314_/Q _13174_/A _13722_/B1 _13519_/X _13525_/X vssd1 vssd1 vccd1 vccd1
+ _13526_/Y sky130_fd_sc_hd__a2111oi_2
X_10738_ _18897_/Q _10816_/A2 _12766_/A0 vssd1 vssd1 vccd1 vccd1 _10738_/X sky130_fd_sc_hd__o21a_1
X_17294_ _17292_/Y _17293_/X _17198_/A vssd1 vssd1 vccd1 vccd1 _19448_/D sky130_fd_sc_hd__a21oi_1
XFILLER_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19033_ _19647_/CLK _19033_/D vssd1 vssd1 vccd1 vccd1 _19033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13457_ _19312_/Q _13754_/A2 _13722_/B1 _13450_/X _13456_/X vssd1 vssd1 vccd1 vccd1
+ _13457_/Y sky130_fd_sc_hd__a2111oi_2
X_16245_ _17676_/A0 _18860_/Q _16245_/S vssd1 vssd1 vccd1 vccd1 _18860_/D sky130_fd_sc_hd__mux2_1
X_10669_ _11601_/A _10669_/B vssd1 vssd1 vccd1 vccd1 _10669_/Y sky130_fd_sc_hd__nor2_1
X_12408_ _12408_/A _12408_/B vssd1 vssd1 vccd1 vccd1 _12408_/X sky130_fd_sc_hd__or2_1
X_16176_ _17706_/A0 _18793_/Q _16193_/S vssd1 vssd1 vccd1 vccd1 _18793_/D sky130_fd_sc_hd__mux2_1
X_13388_ _13312_/A _14146_/A _13909_/B1 vssd1 vssd1 vccd1 vccd1 _13388_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12339_ _18373_/Q _12432_/B1 _09992_/B _08858_/A vssd1 vssd1 vccd1 vccd1 _12340_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_5_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15127_ _14224_/B _12312_/X _16156_/B vssd1 vssd1 vccd1 vccd1 _15127_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15058_ _18542_/Q _17669_/A0 _15078_/S vssd1 vssd1 vccd1 vccd1 _18542_/D sky130_fd_sc_hd__mux2_1
XFILLER_269_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _17969_/Q _14036_/A _14008_/Y _14037_/C1 vssd1 vssd1 vccd1 vccd1 _17969_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_268_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18817_ _18817_/CLK _18817_/D vssd1 vssd1 vccd1 vccd1 _18817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09550_ _18445_/Q _18346_/Q _11160_/S vssd1 vssd1 vccd1 vccd1 _09550_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18748_ _18749_/CLK _18748_/D vssd1 vssd1 vccd1 vccd1 _18748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_283_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09481_ _09992_/A _09481_/B vssd1 vssd1 vccd1 vccd1 _09481_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18679_ _18683_/CLK _18679_/D vssd1 vssd1 vccd1 vccd1 _18679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1309 _11972_/X vssd1 vssd1 vccd1 vccd1 _15881_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09817_ _13263_/A _09818_/B vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__nand2_2
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09748_ _18239_/Q _18814_/Q _09770_/S vssd1 vssd1 vccd1 vccd1 _09748_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09679_ _11161_/S _09674_/X _09678_/X vssd1 vssd1 vccd1 vccd1 _09679_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_95_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _17982_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11710_ _18531_/Q _18530_/Q vssd1 vssd1 vccd1 vccd1 _11711_/B sky130_fd_sc_hd__nand2_2
XFILLER_55_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12603_/B _11626_/Y _13911_/A vssd1 vssd1 vccd1 vccd1 _12690_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19099_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_202_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11641_ _13761_/A vssd1 vssd1 vccd1 vccd1 _11641_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_199_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14360_ _18212_/Q _16501_/A0 _14382_/S vssd1 vssd1 vccd1 vccd1 _18212_/D sky130_fd_sc_hd__mux2_1
X_11572_ _11572_/A1 _18164_/Q _18810_/Q _10856_/C _11584_/C1 vssd1 vssd1 vccd1 vccd1
+ _11572_/X sky130_fd_sc_hd__a221o_1
XFILLER_211_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13311_ _13311_/A _13311_/B vssd1 vssd1 vccd1 vccd1 _14144_/B sky130_fd_sc_hd__xnor2_1
XFILLER_182_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10523_ _11365_/B2 _16617_/A0 _10522_/X _11133_/B2 vssd1 vssd1 vccd1 vccd1 _13743_/A
+ sky130_fd_sc_hd__o2bb2a_2
Xinput19 core_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14291_ _17709_/A0 _18150_/Q _14305_/S vssd1 vssd1 vccd1 vccd1 _18150_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16030_ _16020_/A _16056_/B _18729_/Q vssd1 vssd1 vccd1 vccd1 _16030_/X sky130_fd_sc_hd__a21o_1
X_13242_ _19532_/Q _13372_/S vssd1 vssd1 vccd1 vccd1 _13242_/X sky130_fd_sc_hd__or2_1
X_10454_ _13797_/S _10454_/B vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__or2_4
XFILLER_136_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13173_ _19368_/Q _13247_/A2 _13171_/X _13172_/X _13247_/C1 vssd1 vssd1 vccd1 vccd1
+ _13174_/C sky130_fd_sc_hd__o221a_2
X_10385_ _17946_/Q _11451_/A2 _10384_/X vssd1 vssd1 vccd1 vccd1 _10385_/X sky130_fd_sc_hd__o21a_4
XFILLER_184_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12124_ _17835_/Q _12122_/B _12123_/Y vssd1 vssd1 vccd1 vccd1 _17835_/D sky130_fd_sc_hd__o21a_1
XFILLER_124_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17981_ _17982_/CLK _17981_/D vssd1 vssd1 vccd1 vccd1 _17981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16932_ _17346_/A _16932_/B vssd1 vssd1 vccd1 vccd1 _19317_/D sky130_fd_sc_hd__and2_1
Xfanout1810 _17380_/A vssd1 vssd1 vccd1 vccd1 _17376_/A sky130_fd_sc_hd__buf_4
X_12055_ _17805_/Q _12085_/B vssd1 vssd1 vccd1 vccd1 _12055_/X sky130_fd_sc_hd__or2_1
Xfanout1821 _14340_/A vssd1 vssd1 vccd1 vccd1 _13100_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1832 _17336_/A vssd1 vssd1 vccd1 vccd1 _17326_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1843 _13987_/C1 vssd1 vssd1 vccd1 vccd1 _12428_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11006_ _11004_/X _11005_/X _11478_/S vssd1 vssd1 vccd1 vccd1 _11006_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1854 _13987_/C1 vssd1 vssd1 vccd1 vccd1 _16960_/A sky130_fd_sc_hd__buf_4
Xfanout1865 _16812_/B1 vssd1 vssd1 vccd1 vccd1 _16964_/A sky130_fd_sc_hd__buf_4
X_16863_ _16892_/A _16863_/B vssd1 vssd1 vccd1 vccd1 _19300_/D sky130_fd_sc_hd__and2_1
XFILLER_238_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1876 _14423_/B vssd1 vssd1 vccd1 vccd1 _17261_/A sky130_fd_sc_hd__buf_4
XFILLER_238_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1887 _16142_/B1 vssd1 vssd1 vccd1 vccd1 _16149_/A sky130_fd_sc_hd__buf_4
Xfanout1898 _16740_/A vssd1 vssd1 vccd1 vccd1 _16752_/A sky130_fd_sc_hd__buf_4
XFILLER_237_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18602_ _19047_/CLK _18602_/D vssd1 vssd1 vccd1 vccd1 _18602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15814_ _18606_/Q _17704_/A0 _15832_/S vssd1 vssd1 vccd1 vccd1 _18606_/D sky130_fd_sc_hd__mux2_1
XFILLER_219_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19582_ _19614_/CLK _19582_/D vssd1 vssd1 vccd1 vccd1 _19582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16794_ _19286_/Q _16794_/B vssd1 vssd1 vccd1 vccd1 _16799_/C sky130_fd_sc_hd__and2_2
XFILLER_253_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18533_ _19047_/CLK _18533_/D vssd1 vssd1 vccd1 vccd1 _18533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_218_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _15728_/A _15728_/B _15723_/B vssd1 vssd1 vccd1 vccd1 _15749_/B sky130_fd_sc_hd__o21ba_1
XFILLER_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _12957_/A _12957_/B vssd1 vssd1 vccd1 vccd1 _14141_/D sky130_fd_sc_hd__xor2_4
XFILLER_206_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18464_ _19643_/CLK _18464_/D vssd1 vssd1 vccd1 vccd1 _18464_/Q sky130_fd_sc_hd__dfxtp_1
X_11908_ _11908_/A _11908_/B vssd1 vssd1 vccd1 vccd1 _11909_/B sky130_fd_sc_hd__nor2_8
XFILLER_233_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15676_ _18587_/Q _15800_/A2 _15675_/X _15718_/C1 vssd1 vssd1 vccd1 vccd1 _18587_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12888_ _12888_/A vssd1 vssd1 vccd1 vccd1 _12888_/Y sky130_fd_sc_hd__inv_2
XANTENNA_260 input217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_271 input235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_282 input244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17415_ _11740_/Y _15118_/A _15117_/A _17795_/Q _15116_/B vssd1 vssd1 vccd1 vccd1
+ _17415_/X sky130_fd_sc_hd__a221o_1
X_14627_ _17686_/A0 _18434_/Q _14630_/S vssd1 vssd1 vccd1 vccd1 _18434_/D sky130_fd_sc_hd__mux2_1
XFILLER_221_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_293 _11950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11839_ _11887_/B1 _11837_/X _11838_/X vssd1 vssd1 vccd1 vccd1 _11840_/B sky130_fd_sc_hd__a21oi_4
X_18395_ _19399_/CLK _18395_/D vssd1 vssd1 vccd1 vccd1 _18395_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17346_ _17346_/A _17346_/B vssd1 vssd1 vccd1 vccd1 _19470_/D sky130_fd_sc_hd__and2_1
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14558_ _14592_/A _14558_/B vssd1 vssd1 vccd1 vccd1 _18387_/D sky130_fd_sc_hd__or2_1
XFILLER_174_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13509_ _13322_/Y _13491_/Y _13508_/X _13490_/X _13968_/B2 vssd1 vssd1 vccd1 vccd1
+ _13509_/X sky130_fd_sc_hd__a32o_1
XFILLER_186_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17277_ _19443_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17277_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14489_ _16393_/A _17691_/B vssd1 vssd1 vccd1 vccd1 _14489_/Y sky130_fd_sc_hd__nand2_2
X_19016_ _19208_/CLK _19016_/D vssd1 vssd1 vccd1 vccd1 _19016_/Q sky130_fd_sc_hd__dfxtp_1
X_16228_ _16592_/A0 _18843_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _18843_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16159_ _15416_/A _15116_/A _16156_/Y _16158_/X vssd1 vssd1 vccd1 vccd1 _16159_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08981_ _11513_/A1 _18605_/Q _18176_/Q _11503_/S0 vssd1 vssd1 vccd1 vccd1 _08981_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09602_ _19072_/Q _18976_/Q _10717_/S vssd1 vssd1 vccd1 vccd1 _09602_/X sky130_fd_sc_hd__mux2_1
XFILLER_272_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09533_ _11157_/A1 _19137_/Q _11160_/S _19105_/Q vssd1 vssd1 vccd1 vccd1 _09533_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_260_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09464_ _18850_/Q _18882_/Q _09464_/S vssd1 vssd1 vccd1 vccd1 _09464_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09395_ _10346_/S _09388_/X _09387_/X _10356_/C1 vssd1 vssd1 vccd1 vccd1 _09395_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_269_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_142_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19650_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_279_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10170_ _19064_/Q _19032_/Q _10176_/S vssd1 vssd1 vccd1 vccd1 _10170_/X sky130_fd_sc_hd__mux2_1
Xoutput470 _18129_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[28] sky130_fd_sc_hd__buf_4
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput481 _18110_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[9] sky130_fd_sc_hd__buf_4
Xfanout1106 _12588_/Y vssd1 vssd1 vccd1 vccd1 _13930_/B1 sky130_fd_sc_hd__buf_6
XFILLER_133_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1117 _12451_/X vssd1 vssd1 vccd1 vccd1 _13941_/B sky130_fd_sc_hd__buf_4
XFILLER_266_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1128 _15124_/B vssd1 vssd1 vccd1 vccd1 _15140_/B sky130_fd_sc_hd__clkbuf_4
Xfanout1139 _09437_/B vssd1 vssd1 vccd1 vccd1 _16500_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_259_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13860_ _13860_/A _13860_/B vssd1 vssd1 vccd1 vccd1 _14150_/B sky130_fd_sc_hd__xor2_2
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12811_ _12748_/A _12810_/Y _12935_/S vssd1 vssd1 vccd1 vccd1 _12811_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13791_ _13791_/A _13791_/B _13791_/C vssd1 vssd1 vccd1 vccd1 _13791_/X sky130_fd_sc_hd__and3_1
XFILLER_90_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _15531_/A _15531_/B vssd1 vssd1 vccd1 vccd1 _15530_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12445_/B _12740_/X _09075_/X vssd1 vssd1 vccd1 vccd1 _13483_/B sky130_fd_sc_hd__a21o_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12600_/B _12639_/B _12729_/B vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__mux2_1
X_15461_ _15268_/B _15365_/X _15457_/Y _15458_/Y _15460_/Y vssd1 vssd1 vccd1 vccd1
+ _15558_/A sky130_fd_sc_hd__a311oi_4
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17200_ _19418_/Q fanout533/X _17199_/Y _17119_/B vssd1 vssd1 vccd1 vccd1 _17201_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14412_ _16619_/A0 _18263_/Q _14412_/S vssd1 vssd1 vccd1 vccd1 _18263_/D sky130_fd_sc_hd__mux2_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11624_/A1 _17723_/A0 _11623_/X _09523_/A vssd1 vssd1 vccd1 vccd1 _13941_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_169_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18180_ _19589_/CLK _18180_/D vssd1 vssd1 vccd1 vccd1 _18180_/Q sky130_fd_sc_hd__dfxtp_1
X_15392_ _12788_/B _15391_/Y _15437_/B1 vssd1 vssd1 vccd1 vccd1 _15392_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_129_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17131_ _17559_/B _17120_/Y _17130_/Y _17231_/A vssd1 vssd1 vccd1 vccd1 _17131_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11555_ _13908_/A _11555_/B vssd1 vssd1 vccd1 vccd1 _13938_/B sky130_fd_sc_hd__xnor2_4
X_14343_ _15039_/A _14345_/B _14343_/C vssd1 vssd1 vccd1 vccd1 _18198_/D sky130_fd_sc_hd__and3_4
XFILLER_183_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10506_ _18261_/Q _18836_/Q _10511_/S vssd1 vssd1 vccd1 vccd1 _10506_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17062_ _17567_/A _17074_/A2 _17061_/X _17322_/A vssd1 vssd1 vccd1 vccd1 _19364_/D
+ sky130_fd_sc_hd__o211a_1
X_14274_ _16592_/A0 _18133_/Q _14277_/S vssd1 vssd1 vccd1 vccd1 _18133_/D sky130_fd_sc_hd__mux2_1
X_11486_ _10009_/A _11475_/X _11483_/Y _11485_/Y vssd1 vssd1 vccd1 vccd1 _11486_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16013_ _18722_/Q _16019_/A2 _16012_/X _14197_/A vssd1 vssd1 vccd1 vccd1 _18722_/D
+ sky130_fd_sc_hd__o211a_1
X_13225_ _13225_/A _13225_/B _13225_/C vssd1 vssd1 vccd1 vccd1 _13226_/B sky130_fd_sc_hd__or3_1
XFILLER_170_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10437_ _18869_/Q _18901_/Q _11598_/S vssd1 vssd1 vccd1 vccd1 _10437_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ _13136_/S _13135_/X _13197_/B1 vssd1 vssd1 vccd1 vccd1 _13156_/Y sky130_fd_sc_hd__o21bai_2
X_10368_ _10373_/S _10363_/X _10367_/X _08895_/A vssd1 vssd1 vccd1 vccd1 _10368_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12107_ _12107_/A _12112_/C vssd1 vssd1 vccd1 vccd1 _12107_/Y sky130_fd_sc_hd__nor2_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17964_ _18627_/CLK _17964_/D vssd1 vssd1 vccd1 vccd1 _17964_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _12873_/Y _12877_/Y _13130_/A vssd1 vssd1 vccd1 vccd1 _13087_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10299_ _19646_/Q _18935_/Q _10299_/S vssd1 vssd1 vccd1 vccd1 _10299_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16915_ _19313_/Q _17172_/B _16967_/S vssd1 vssd1 vccd1 vccd1 _16916_/B sky130_fd_sc_hd__mux2_1
Xfanout1640 _08857_/Y vssd1 vssd1 vccd1 vccd1 _09012_/A sky130_fd_sc_hd__clkbuf_4
X_12038_ _17894_/Q _12035_/B _12037_/X _12383_/C1 vssd1 vssd1 vccd1 vccd1 _17796_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1651 _10366_/A1 vssd1 vssd1 vccd1 vccd1 _10294_/A1 sky130_fd_sc_hd__buf_6
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17895_ _17901_/CLK _17895_/D vssd1 vssd1 vccd1 vccd1 _17895_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1662 _08850_/Y vssd1 vssd1 vccd1 vccd1 _09873_/A1 sky130_fd_sc_hd__buf_12
Xfanout1673 _11607_/S vssd1 vssd1 vccd1 vccd1 _10746_/S sky130_fd_sc_hd__buf_12
XFILLER_265_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1684 _10625_/A1 vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__buf_12
X_19634_ _19634_/CLK _19634_/D vssd1 vssd1 vccd1 vccd1 _19634_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1695 _08845_/Y vssd1 vssd1 vccd1 vccd1 _11404_/A1 sky130_fd_sc_hd__buf_6
X_16846_ _16967_/S _16846_/B vssd1 vssd1 vccd1 vccd1 _16846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19565_ _19565_/CLK _19565_/D vssd1 vssd1 vccd1 vccd1 _19565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16777_ _19280_/Q _16778_/B vssd1 vssd1 vccd1 vccd1 _16779_/B sky130_fd_sc_hd__nor2_1
XFILLER_253_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13989_ _17959_/Q _14020_/B _13988_/Y _14037_/C1 vssd1 vssd1 vccd1 vccd1 _17959_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18516_ _18517_/CLK _18516_/D vssd1 vssd1 vccd1 vccd1 _18516_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15728_ _15728_/A _15728_/B vssd1 vssd1 vccd1 vccd1 _15728_/Y sky130_fd_sc_hd__xnor2_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19496_ _19534_/CLK _19496_/D vssd1 vssd1 vccd1 vccd1 _19496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18447_ _19594_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15659_ _15744_/A _15687_/B vssd1 vssd1 vccd1 vccd1 _15686_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09180_ _18058_/Q _10101_/B _09179_/X _10335_/S vssd1 vssd1 vccd1 vccd1 _09180_/X
+ sky130_fd_sc_hd__o211a_1
X_18378_ _19483_/CLK _18378_/D vssd1 vssd1 vccd1 vccd1 _18378_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_187_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17329_ _08818_/Y _16870_/Y _17377_/S vssd1 vssd1 vccd1 vccd1 _17330_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_1__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_1__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08964_ _11511_/A _08959_/X _08963_/X vssd1 vssd1 vccd1 vccd1 _08964_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_248_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput209 localMemory_wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08895_ _08895_/A _12023_/A vssd1 vssd1 vccd1 vccd1 _08895_/Y sky130_fd_sc_hd__nor2_2
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09516_ _09723_/S _09515_/X _09514_/X _09978_/A1 vssd1 vssd1 vccd1 vccd1 _09516_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_25_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09447_ _18023_/Q _17991_/Q _09464_/S vssd1 vssd1 vccd1 vccd1 _09447_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ _10297_/A1 _09368_/X _09369_/X vssd1 vssd1 vccd1 vccd1 _09378_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11340_ _11360_/A1 _18321_/Q _17772_/Q _11340_/B2 vssd1 vssd1 vccd1 vccd1 _11340_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11271_ _18858_/Q _18890_/Q _19050_/Q _19018_/Q _11284_/B2 _11622_/A1 vssd1 vssd1
+ vccd1 vccd1 _11271_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _15905_/A _12536_/Y _12505_/Y vssd1 vssd1 vccd1 vccd1 _13010_/X sky130_fd_sc_hd__a21o_1
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10222_ _10297_/A1 _10212_/X _10213_/X vssd1 vssd1 vccd1 vccd1 _10222_/X sky130_fd_sc_hd__o21a_1
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10153_ _10747_/A1 _10152_/X _11501_/B1 vssd1 vssd1 vccd1 vccd1 _10153_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14961_ _18497_/Q _15011_/A2 _14960_/Y _16787_/A vssd1 vssd1 vccd1 vccd1 _18497_/D
+ sky130_fd_sc_hd__a211o_1
X_10084_ _11218_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__nor2_1
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16700_ _19252_/Q _16697_/B _16698_/Y vssd1 vssd1 vccd1 vccd1 _19252_/D sky130_fd_sc_hd__o21a_1
XFILLER_236_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13912_ _10160_/A _13912_/A2 _13912_/B1 vssd1 vssd1 vccd1 vccd1 _13913_/B sky130_fd_sc_hd__a21oi_1
XFILLER_208_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17680_ _17680_/A0 _19607_/Q _17690_/S vssd1 vssd1 vccd1 vccd1 _19607_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14892_ _17810_/Q _15002_/B _14891_/X vssd1 vssd1 vccd1 vccd1 _14892_/X sky130_fd_sc_hd__o21a_1
XFILLER_262_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16631_ _17724_/A _19232_/Q _16630_/Y vssd1 vssd1 vccd1 vccd1 _19232_/D sky130_fd_sc_hd__o21a_1
XFILLER_235_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13843_ _13843_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _13843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19350_ _19483_/CLK _19350_/D vssd1 vssd1 vccd1 vccd1 _19350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16562_ _17695_/A0 _19166_/Q _16590_/S vssd1 vssd1 vccd1 vccd1 _19166_/D sky130_fd_sc_hd__mux2_1
X_10986_ _09574_/A _09151_/X _11143_/A1 vssd1 vssd1 vccd1 vccd1 _10988_/A sky130_fd_sc_hd__a21oi_1
X_13774_ _17945_/Q _13940_/A2 _13773_/X _14179_/A vssd1 vssd1 vccd1 vccd1 _17945_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18301_ _19453_/CLK _18301_/D vssd1 vssd1 vccd1 vccd1 _18301_/Q sky130_fd_sc_hd__dfxtp_1
X_15513_ _18579_/Q _15512_/C _18580_/Q vssd1 vssd1 vccd1 vccd1 _15514_/B sky130_fd_sc_hd__a21oi_1
XFILLER_71_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19281_ _19285_/CLK _19281_/D vssd1 vssd1 vccd1 vccd1 _19281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12725_ _12823_/B _12723_/X _12823_/A vssd1 vssd1 vccd1 vccd1 _12726_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16493_ _16526_/A0 _19099_/Q _16515_/S vssd1 vssd1 vccd1 vccd1 _19099_/D sky130_fd_sc_hd__mux2_1
X_18232_ _19159_/CLK _18232_/D vssd1 vssd1 vccd1 vccd1 _18232_/Q sky130_fd_sc_hd__dfxtp_1
X_15444_ _15444_/A _15444_/B vssd1 vssd1 vccd1 vccd1 _15445_/B sky130_fd_sc_hd__nand2_1
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12656_ _12656_/A _12656_/B _13891_/A _13860_/A vssd1 vssd1 vccd1 vccd1 _12656_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_90_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18163_ _19628_/CLK _18163_/D vssd1 vssd1 vccd1 vccd1 _18163_/Q sky130_fd_sc_hd__dfxtp_1
X_11607_ _11603_/X _11606_/X _11607_/S vssd1 vssd1 vccd1 vccd1 _11607_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12587_ _12756_/B _12587_/B vssd1 vssd1 vccd1 vccd1 _12587_/Y sky130_fd_sc_hd__nand2_2
X_15375_ _19467_/Q _19401_/Q _15374_/X vssd1 vssd1 vccd1 vccd1 _15376_/B sky130_fd_sc_hd__o21ai_4
XFILLER_168_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17114_ _17211_/B _17114_/A2 _17113_/X _17322_/A vssd1 vssd1 vccd1 vccd1 _19390_/D
+ sky130_fd_sc_hd__o211a_1
X_14326_ _18183_/Q _17710_/A0 _14338_/S vssd1 vssd1 vccd1 vccd1 _18183_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18094_ _19306_/CLK _18094_/D vssd1 vssd1 vccd1 vccd1 _18094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11538_ _13597_/A _11673_/B _11534_/B _13616_/A _11536_/X vssd1 vssd1 vccd1 vccd1
+ _11669_/B sky130_fd_sc_hd__a41o_4
XFILLER_117_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17045_ _19359_/Q _17045_/B vssd1 vssd1 vccd1 vccd1 _17045_/X sky130_fd_sc_hd__or2_1
X_11469_ _11469_/A1 _19630_/Q _18919_/Q _11477_/S vssd1 vssd1 vccd1 vccd1 _11470_/B
+ sky130_fd_sc_hd__a22o_1
X_14257_ _18300_/Q _14261_/A2 _14256_/X _14450_/B vssd1 vssd1 vccd1 vccd1 _18126_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13208_ _19531_/Q _13921_/S vssd1 vssd1 vccd1 vccd1 _13208_/X sky130_fd_sc_hd__or2_1
XFILLER_125_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14188_ _18705_/Q _18092_/Q _14200_/S vssd1 vssd1 vccd1 vccd1 _14189_/B sky130_fd_sc_hd__mux2_1
XFILLER_140_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _13139_/A vssd1 vssd1 vccd1 vccd1 _13139_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ _19092_/CLK _18996_/D vssd1 vssd1 vccd1 vccd1 _18996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17947_ _18627_/CLK _17947_/D vssd1 vssd1 vccd1 vccd1 _17947_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1470 _10656_/S vssd1 vssd1 vccd1 vccd1 _10667_/S sky130_fd_sc_hd__buf_6
XFILLER_39_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1481 fanout1485/X vssd1 vssd1 vccd1 vccd1 _11284_/B2 sky130_fd_sc_hd__buf_6
X_17878_ _19320_/CLK _17878_/D vssd1 vssd1 vccd1 vccd1 _17878_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1492 _10721_/S vssd1 vssd1 vccd1 vccd1 _10717_/S sky130_fd_sc_hd__buf_6
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16829_ _16821_/A _17819_/Q _12476_/Y vssd1 vssd1 vccd1 vccd1 _16831_/A sky130_fd_sc_hd__a21o_1
X_19617_ _19618_/CLK _19617_/D vssd1 vssd1 vccd1 vccd1 _19617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19548_ _19553_/CLK _19548_/D vssd1 vssd1 vccd1 vccd1 _19548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ _11498_/A1 _19563_/Q _09306_/S _19595_/Q _09374_/S vssd1 vssd1 vccd1 vccd1
+ _09301_/X sky130_fd_sc_hd__o221a_1
XFILLER_206_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19479_ _19481_/CLK _19479_/D vssd1 vssd1 vccd1 vccd1 _19479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09232_ _09232_/A _09232_/B vssd1 vssd1 vccd1 vccd1 _09232_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09163_ _09161_/X _09162_/X _10169_/S vssd1 vssd1 vccd1 vccd1 _09163_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09094_ _14074_/C _09542_/S vssd1 vssd1 vccd1 vccd1 _09094_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_147_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09996_ _10027_/A _18016_/Q vssd1 vssd1 vccd1 vccd1 _09996_/X sky130_fd_sc_hd__or2_1
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _08947_/A _08947_/B vssd1 vssd1 vccd1 vccd1 _08947_/X sky130_fd_sc_hd__or2_4
XFILLER_88_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ _15549_/A _12442_/A vssd1 vssd1 vccd1 vccd1 _12320_/C sky130_fd_sc_hd__or2_2
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10840_ _18646_/Q _18068_/Q _10840_/S vssd1 vssd1 vccd1 vccd1 _10840_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10771_ _18864_/Q _18896_/Q _10856_/C vssd1 vssd1 vccd1 vccd1 _10771_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12510_ _12548_/A _12575_/A vssd1 vssd1 vccd1 vccd1 _12510_/X sky130_fd_sc_hd__or2_4
XFILLER_197_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13490_ _13483_/Y _13486_/Y _13489_/X _13966_/C1 vssd1 vssd1 vccd1 vccd1 _13490_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12441_ _12756_/A _12455_/A vssd1 vssd1 vccd1 vccd1 _12441_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12372_ _18384_/Q _12420_/B1 _09046_/B _18201_/Q vssd1 vssd1 vccd1 vccd1 _12373_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_15160_ _15149_/Y _15156_/X _15159_/Y vssd1 vssd1 vccd1 vccd1 _15163_/A sky130_fd_sc_hd__o21a_1
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14111_ _16594_/A0 _18050_/Q _14131_/S vssd1 vssd1 vccd1 vccd1 _18050_/D sky130_fd_sc_hd__mux2_1
X_11323_ _18608_/Q _18179_/Q _11325_/S vssd1 vssd1 vccd1 vccd1 _11323_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15091_ _19386_/Q _15092_/B _15091_/C vssd1 vssd1 vccd1 vccd1 _15093_/D sky130_fd_sc_hd__and3_2
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11254_ _11234_/X _11237_/X _11253_/X vssd1 vssd1 vccd1 vccd1 _11254_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14042_ _16526_/A0 _17984_/Q _14064_/S vssd1 vssd1 vccd1 vccd1 _17984_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10205_ _10203_/X _10204_/X _10205_/S vssd1 vssd1 vccd1 vccd1 _10205_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18850_ _19614_/CLK _18850_/D vssd1 vssd1 vccd1 vccd1 _18850_/Q sky130_fd_sc_hd__dfxtp_1
X_11185_ _11190_/A1 _18610_/Q _18181_/Q _09883_/B vssd1 vssd1 vccd1 vccd1 _11185_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_267_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17801_ _18201_/CLK _17801_/D vssd1 vssd1 vccd1 vccd1 _17801_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_268_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10136_ _11046_/S1 _10125_/X _10135_/X _11438_/B1 vssd1 vssd1 vccd1 vccd1 _10136_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18781_ _19197_/CLK _18781_/D vssd1 vssd1 vccd1 vccd1 _18781_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15993_ _18712_/Q _16005_/A2 _15992_/X _14205_/A vssd1 vssd1 vccd1 vccd1 _18712_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ _18632_/Q vssd1 vssd1 vccd1 vccd1 _18632_/D sky130_fd_sc_hd__clkbuf_2
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10067_ _14141_/A _11651_/B _09897_/Y _12838_/S vssd1 vssd1 vccd1 vccd1 _10068_/B
+ sky130_fd_sc_hd__a211o_1
X_14944_ _14942_/X _14943_/X _14714_/B vssd1 vssd1 vccd1 vccd1 _14944_/X sky130_fd_sc_hd__a21o_1
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17663_ _17663_/A0 _19590_/Q _17687_/S vssd1 vssd1 vccd1 vccd1 _19590_/D sky130_fd_sc_hd__mux2_1
XFILLER_263_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14875_ _14875_/A1 _14874_/X _14875_/B1 vssd1 vssd1 vccd1 vccd1 _14875_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19402_ _19530_/CLK _19402_/D vssd1 vssd1 vccd1 vccd1 _19402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16614_ _16614_/A0 _19217_/Q _16619_/S vssd1 vssd1 vccd1 vccd1 _19217_/D sky130_fd_sc_hd__mux2_1
X_13826_ _19451_/Q _13949_/A2 _13824_/X _13825_/X _13949_/C1 vssd1 vssd1 vccd1 vccd1
+ _13826_/X sky130_fd_sc_hd__o221a_2
X_17594_ _19538_/Q _17622_/A2 _17591_/X _17169_/B _17593_/X vssd1 vssd1 vccd1 vccd1
+ _19538_/D sky130_fd_sc_hd__o221a_1
XFILLER_251_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19333_ _19534_/CLK _19333_/D vssd1 vssd1 vccd1 vccd1 _19333_/Q sky130_fd_sc_hd__dfxtp_1
X_16545_ _16545_/A0 _19150_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _19150_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ _13757_/A _14024_/B vssd1 vssd1 vccd1 vccd1 _13757_/X sky130_fd_sc_hd__or2_4
X_10969_ _11355_/A1 _10966_/X _10968_/X vssd1 vssd1 vccd1 vccd1 _10977_/B sky130_fd_sc_hd__a21oi_1
XFILLER_204_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19264_ _19268_/CLK _19264_/D vssd1 vssd1 vccd1 vccd1 _19264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12708_ _09984_/B _12660_/B _12835_/A vssd1 vssd1 vccd1 vccd1 _12708_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16476_ _16476_/A0 _19083_/Q _16485_/S vssd1 vssd1 vccd1 vccd1 _19083_/D sky130_fd_sc_hd__mux2_1
X_13688_ _19351_/Q _13883_/A2 _13883_/B1 _19479_/Q _13883_/C1 vssd1 vssd1 vccd1 vccd1
+ _13688_/X sky130_fd_sc_hd__a221o_1
X_18215_ _18543_/CLK _18215_/D vssd1 vssd1 vccd1 vccd1 _18215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15427_ _15404_/B _13408_/Y _15133_/B _15426_/X vssd1 vssd1 vccd1 vccd1 _15427_/X
+ sky130_fd_sc_hd__a31o_1
X_12639_ _10753_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _12639_/Y sky130_fd_sc_hd__nand2b_2
X_19195_ _19195_/CLK _19195_/D vssd1 vssd1 vccd1 vccd1 _19195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18146_ _19208_/CLK _18146_/D vssd1 vssd1 vccd1 vccd1 _18146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15358_ _15404_/B _13327_/X _15381_/A3 _15357_/Y vssd1 vssd1 vccd1 vccd1 _15358_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_129_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14309_ _18166_/Q _17693_/A0 _14335_/S vssd1 vssd1 vccd1 vccd1 _18166_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18077_ _19613_/CLK _18077_/D vssd1 vssd1 vccd1 vccd1 _18077_/Q sky130_fd_sc_hd__dfxtp_1
X_15289_ _15289_/A _15289_/B vssd1 vssd1 vccd1 vccd1 _15310_/A sky130_fd_sc_hd__or2_1
XFILLER_132_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17028_ _17187_/B _17032_/A2 _17027_/X _17592_/B vssd1 vssd1 vccd1 vccd1 _19350_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout707 _12543_/X vssd1 vssd1 vccd1 vccd1 _13944_/B sky130_fd_sc_hd__buf_6
X_09850_ _18534_/Q _18409_/Q _10001_/S vssd1 vssd1 vccd1 vccd1 _09850_/X sky130_fd_sc_hd__mux2_1
Xfanout718 _13952_/A2 vssd1 vssd1 vccd1 vccd1 _13754_/A2 sky130_fd_sc_hd__buf_4
Xfanout729 _16538_/A0 vssd1 vssd1 vccd1 vccd1 _17671_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_259_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09781_ _11284_/A1 _19198_/Q _19166_/Q _09797_/S _10030_/C1 vssd1 vssd1 vccd1 vccd1
+ _09781_/X sky130_fd_sc_hd__a221o_1
X_18979_ _19075_/CLK _18979_/D vssd1 vssd1 vccd1 vccd1 _18979_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09215_ _18636_/Q _18058_/Q _10353_/S vssd1 vssd1 vccd1 vccd1 _09215_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09146_ input125/X input160/X _09657_/S vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__mux2_8
XFILLER_154_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09077_ _12455_/A _12740_/C _12740_/A vssd1 vssd1 vccd1 vccd1 _12445_/A sky130_fd_sc_hd__a21o_4
XFILLER_146_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_49_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19614_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09979_ _11495_/B1 _09977_/X _09978_/X _09958_/X _09964_/X vssd1 vssd1 vccd1 vccd1
+ _09979_/X sky130_fd_sc_hd__o32a_4
XFILLER_264_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12990_ _13314_/S _12990_/B vssd1 vssd1 vccd1 vccd1 _12990_/X sky130_fd_sc_hd__or2_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11941_ _14667_/A1 _11863_/B _11863_/C _11953_/A2 input228/X vssd1 vssd1 vccd1 vccd1
+ _11941_/X sky130_fd_sc_hd__a32o_4
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _16619_/A0 _18466_/Q _14660_/S vssd1 vssd1 vccd1 vccd1 _18466_/D sky130_fd_sc_hd__mux2_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11872_ _11909_/A _11872_/B vssd1 vssd1 vccd1 vccd1 _11872_/X sky130_fd_sc_hd__and2_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _13904_/A _13611_/B vssd1 vssd1 vccd1 vccd1 _13611_/X sky130_fd_sc_hd__or2_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ _10663_/S _10812_/X _10813_/X vssd1 vssd1 vccd1 vccd1 _10823_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14591_ _18404_/Q _14591_/A2 _14591_/B1 input34/X vssd1 vssd1 vccd1 vccd1 _14592_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16330_ _18942_/Q _16529_/A0 _16358_/S vssd1 vssd1 vccd1 vccd1 _18942_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13542_ _13606_/C _13542_/B vssd1 vssd1 vccd1 vccd1 _13542_/X sky130_fd_sc_hd__or2_1
X_10754_ _10754_/A _10754_/B vssd1 vssd1 vccd1 vccd1 _12638_/A sky130_fd_sc_hd__nor2_8
XFILLER_213_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16261_ _17692_/A0 _18875_/Q _16292_/S vssd1 vssd1 vccd1 vccd1 _18875_/D sky130_fd_sc_hd__mux2_1
X_13473_ _14238_/A _13479_/C vssd1 vssd1 vccd1 vccd1 _13473_/Y sky130_fd_sc_hd__xnor2_2
X_10685_ _10683_/X _10684_/X _11248_/S vssd1 vssd1 vccd1 vccd1 _10685_/X sky130_fd_sc_hd__mux2_1
X_18000_ _19602_/CLK _18000_/D vssd1 vssd1 vccd1 vccd1 _18000_/Q sky130_fd_sc_hd__dfxtp_1
X_15212_ _18567_/Q _15351_/A2 _15211_/X _14430_/B vssd1 vssd1 vccd1 vccd1 _18567_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12424_ _12427_/A _12424_/B vssd1 vssd1 vccd1 vccd1 _12424_/Y sky130_fd_sc_hd__nand2_1
X_16192_ _16622_/A0 _18809_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _18809_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15143_ _19458_/Q _19392_/Q vssd1 vssd1 vccd1 vccd1 _15167_/A sky130_fd_sc_hd__nand2_1
X_12355_ _12379_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12355_/Y sky130_fd_sc_hd__nand2_1
XFILLER_275_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11306_ _10785_/A _11304_/X _11305_/X _11570_/B1 vssd1 vssd1 vccd1 vccd1 _11306_/X
+ sky130_fd_sc_hd__o31a_1
X_15074_ _18558_/Q _16486_/A0 _15078_/S vssd1 vssd1 vccd1 vccd1 _18558_/D sky130_fd_sc_hd__mux2_1
X_12286_ _18095_/Q _12305_/A2 _12305_/B1 _18518_/Q vssd1 vssd1 vccd1 vccd1 _14681_/C
+ sky130_fd_sc_hd__a22o_4
XFILLER_113_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14025_ _17977_/Q _14028_/A _14024_/Y _14029_/C1 vssd1 vssd1 vccd1 vccd1 _17977_/D
+ sky130_fd_sc_hd__o211a_1
X_18902_ _18902_/CLK _18902_/D vssd1 vssd1 vccd1 vccd1 _18902_/Q sky130_fd_sc_hd__dfxtp_1
X_11237_ _11568_/A _11235_/X _11236_/X _11237_/B1 vssd1 vssd1 vccd1 vccd1 _11237_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11168_ _18252_/Q _11171_/S _09683_/A _11167_/X vssd1 vssd1 vccd1 vccd1 _11168_/X
+ sky130_fd_sc_hd__o211a_1
X_18833_ _19025_/CLK _18833_/D vssd1 vssd1 vccd1 vccd1 _18833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10119_ _11484_/B1 _10097_/X _10105_/Y _10111_/Y _10118_/Y vssd1 vssd1 vccd1 vccd1
+ _10119_/X sky130_fd_sc_hd__a32o_4
X_18764_ _19076_/CLK _18764_/D vssd1 vssd1 vccd1 vccd1 _18764_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ _18703_/Q _15953_/B _15976_/B1 _18752_/Q _15976_/C1 vssd1 vssd1 vccd1 vccd1
+ _15976_/X sky130_fd_sc_hd__a221o_1
X_11099_ _11078_/X _11081_/X _11098_/X vssd1 vssd1 vccd1 vccd1 _11099_/X sky130_fd_sc_hd__a21o_1
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17715_ _17715_/A0 _19641_/Q _17718_/S vssd1 vssd1 vccd1 vccd1 _19641_/D sky130_fd_sc_hd__mux2_1
X_14927_ _14927_/A vssd1 vssd1 vccd1 vccd1 _14927_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_64_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18695_ _18746_/CLK _18695_/D vssd1 vssd1 vccd1 vccd1 _18695_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17646_ _17679_/A0 _19574_/Q _17657_/S vssd1 vssd1 vccd1 vccd1 _19574_/D sky130_fd_sc_hd__mux2_1
XFILLER_282_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14858_ _14696_/A _18271_/Q _14857_/Y _14918_/B1 vssd1 vssd1 vccd1 vccd1 _14858_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_63_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13809_ _17946_/Q _13940_/A2 _13808_/X _14029_/C1 vssd1 vssd1 vccd1 vccd1 _17946_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17577_ _17577_/A _17589_/B vssd1 vssd1 vccd1 vccd1 _17577_/X sky130_fd_sc_hd__or2_1
X_14789_ _17800_/Q _14982_/B vssd1 vssd1 vccd1 vccd1 _14789_/X sky130_fd_sc_hd__or2_1
X_19316_ _19363_/CLK _19316_/D vssd1 vssd1 vccd1 vccd1 _19316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16528_ _16594_/A0 _19133_/Q _16548_/S vssd1 vssd1 vccd1 vccd1 _19133_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19247_ _19280_/CLK _19247_/D vssd1 vssd1 vccd1 vccd1 _19247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16459_ _16459_/A _16459_/B _16459_/C _14074_/B vssd1 vssd1 vccd1 vccd1 _16459_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_192_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09000_ _09043_/A _09031_/S vssd1 vssd1 vccd1 vccd1 _09000_/Y sky130_fd_sc_hd__nor2_2
XFILLER_176_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19178_ _19640_/CLK _19178_/D vssd1 vssd1 vccd1 vccd1 _19178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18129_ _19453_/CLK _18129_/D vssd1 vssd1 vccd1 vccd1 _18129_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_191_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _11556_/B _09902_/B _09902_/C vssd1 vssd1 vccd1 vccd1 _09903_/D sky130_fd_sc_hd__or3_1
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout504 _14667_/A1 vssd1 vssd1 vccd1 vccd1 _11953_/B2 sky130_fd_sc_hd__buf_6
Xfanout515 _17313_/B vssd1 vssd1 vccd1 vccd1 _17289_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_258_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout526 _11769_/B1 vssd1 vssd1 vccd1 vccd1 _11799_/B sky130_fd_sc_hd__buf_4
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout537 _15633_/C1 vssd1 vssd1 vccd1 vccd1 _15782_/B1 sky130_fd_sc_hd__buf_6
X_09833_ _09853_/S _09832_/X _12320_/A vssd1 vssd1 vccd1 vccd1 _09833_/X sky130_fd_sc_hd__a21o_1
XFILLER_141_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout548 _15123_/X vssd1 vssd1 vccd1 vccd1 _15476_/A1 sky130_fd_sc_hd__buf_4
Xfanout559 _15537_/B1 vssd1 vssd1 vccd1 vccd1 _15789_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_274_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09764_ _11568_/A _09764_/B vssd1 vssd1 vccd1 vccd1 _09764_/X sky130_fd_sc_hd__or2_1
XFILLER_100_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_167_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19482_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09695_ _17899_/Q _15120_/A vssd1 vssd1 vccd1 vccd1 _09695_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ _10625_/A1 _18158_/Q _18804_/Q _10619_/S vssd1 vssd1 vccd1 vccd1 _10470_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09129_ _09127_/X _09128_/X _09129_/S vssd1 vssd1 vccd1 vccd1 _09129_/X sky130_fd_sc_hd__mux2_1
X_12140_ _17841_/Q _12138_/B _12139_/Y vssd1 vssd1 vccd1 vccd1 _17841_/D sky130_fd_sc_hd__o21a_1
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12071_ _17813_/Q _12085_/B vssd1 vssd1 vccd1 vccd1 _12071_/X sky130_fd_sc_hd__or2_1
XFILLER_173_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ _09089_/Y _11011_/X _11019_/X _11021_/X vssd1 vssd1 vccd1 vccd1 _11022_/X
+ sky130_fd_sc_hd__o31a_4
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15830_ _18622_/Q _17720_/A0 _15832_/S vssd1 vssd1 vccd1 vccd1 _18622_/D sky130_fd_sc_hd__mux2_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _18591_/Q _15800_/A2 _15760_/X _14449_/B vssd1 vssd1 vccd1 vccd1 _18591_/D
+ sky130_fd_sc_hd__o211a_1
X_12973_ _19364_/Q _13247_/A2 _12971_/X _12972_/X _13247_/C1 vssd1 vssd1 vccd1 vccd1
+ _12973_/X sky130_fd_sc_hd__o221a_4
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _11686_/A _17520_/A2 _17532_/A2 _17812_/Q _17550_/A vssd1 vssd1 vccd1 vccd1
+ _17500_/X sky130_fd_sc_hd__a221o_1
XFILLER_273_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _18628_/Q _14683_/A _14683_/B _14912_/A1 _12865_/Y vssd1 vssd1 vccd1 vccd1
+ _14712_/X sky130_fd_sc_hd__a32o_1
X_18480_ _19321_/CLK _18480_/D vssd1 vssd1 vccd1 vccd1 _18480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _11926_/A1 _11939_/A1 _11820_/B _11935_/B1 input241/X vssd1 vssd1 vccd1 vccd1
+ _11924_/X sky130_fd_sc_hd__a32o_4
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _15672_/A _15672_/B _15671_/A vssd1 vssd1 vccd1 vccd1 _15696_/A sky130_fd_sc_hd__a21oi_2
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_420 _13810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_431 _11849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_442 _13998_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _18570_/Q _17461_/A2 _17546_/A2 vssd1 vssd1 vccd1 vccd1 _17431_/X sky130_fd_sc_hd__o21a_1
X_14643_ _16470_/A0 _18449_/Q _14663_/S vssd1 vssd1 vccd1 vccd1 _18449_/D sky130_fd_sc_hd__mux2_1
XFILLER_221_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_453 _17799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _11859_/B _11819_/X _11794_/Y _11801_/A vssd1 vssd1 vccd1 vccd1 _11855_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_464 _18389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_475 input222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_486 _11929_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10806_ _11112_/A _10804_/X _10805_/X _11361_/S vssd1 vssd1 vccd1 vccd1 _10806_/X
+ sky130_fd_sc_hd__a211o_1
X_17362_ _17592_/B _17362_/B vssd1 vssd1 vccd1 vccd1 _19478_/D sky130_fd_sc_hd__and2_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_497 _14277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14574_ _14576_/A _14574_/B vssd1 vssd1 vccd1 vccd1 _18395_/D sky130_fd_sc_hd__or2_1
XFILLER_242_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11786_ _11820_/A _11807_/B vssd1 vssd1 vccd1 vccd1 _11786_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19101_ _19133_/CLK _19101_/D vssd1 vssd1 vccd1 vccd1 _19101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16313_ _17711_/A0 _18926_/Q _16320_/S vssd1 vssd1 vccd1 vccd1 _18926_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ _19378_/Q _13884_/A2 _13523_/X _13524_/X _13884_/C1 vssd1 vssd1 vccd1 vccd1
+ _13525_/X sky130_fd_sc_hd__o221a_4
X_17293_ _18125_/Q _15717_/B2 _17513_/A _17307_/B vssd1 vssd1 vccd1 vccd1 _17293_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_10737_ _18865_/Q _10744_/S vssd1 vssd1 vccd1 vccd1 _10737_/X sky130_fd_sc_hd__or2_1
XFILLER_158_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19032_ _19647_/CLK _19032_/D vssd1 vssd1 vccd1 vccd1 _19032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16244_ _16608_/A0 _18859_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _18859_/D sky130_fd_sc_hd__mux2_1
X_13456_ _19376_/Q _13951_/A2 _13454_/X _13455_/X _13951_/C1 vssd1 vssd1 vccd1 vccd1
+ _13456_/X sky130_fd_sc_hd__o221a_4
X_10668_ _10666_/X _10667_/X _10668_/S vssd1 vssd1 vccd1 vccd1 _10669_/B sky130_fd_sc_hd__mux2_1
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ _12466_/A0 _12430_/A _12406_/Y _14001_/C1 vssd1 vssd1 vccd1 vccd1 _17910_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16175_ _11376_/B _18792_/Q _16189_/S vssd1 vssd1 vccd1 vccd1 _18792_/D sky130_fd_sc_hd__mux2_1
X_10599_ _13711_/A vssd1 vssd1 vccd1 vccd1 _10599_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13387_ _13387_/A _13387_/B vssd1 vssd1 vccd1 vccd1 _14146_/A sky130_fd_sc_hd__xnor2_1
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15126_ _12312_/X _17211_/A _15731_/B1 _14224_/B vssd1 vssd1 vccd1 vccd1 _15126_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_114_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338_ _17887_/Q _14224_/B vssd1 vssd1 vccd1 vccd1 _12338_/Y sky130_fd_sc_hd__nor2_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15057_ _18541_/Q _16535_/A0 _15078_/S vssd1 vssd1 vccd1 vccd1 _18541_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12269_ _12269_/A _12269_/B _12269_/C input205/X vssd1 vssd1 vccd1 vccd1 _12271_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_269_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14008_ _14036_/A _14008_/B vssd1 vssd1 vccd1 vccd1 _14008_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18816_ _18880_/CLK _18816_/D vssd1 vssd1 vccd1 vccd1 _18816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15959_ _18695_/Q _15977_/A2 _15958_/X _16892_/A vssd1 vssd1 vccd1 vccd1 _18695_/D
+ sky130_fd_sc_hd__o211a_1
X_18747_ _18749_/CLK _18747_/D vssd1 vssd1 vccd1 vccd1 _18747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18678_ _18683_/CLK _18678_/D vssd1 vssd1 vccd1 vccd1 _18678_/Q sky130_fd_sc_hd__dfxtp_1
X_09480_ _09652_/A _09480_/B vssd1 vssd1 vccd1 vccd1 _09481_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17629_ _17662_/A0 _19557_/Q _17648_/S vssd1 vssd1 vccd1 vccd1 _19557_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09816_ _09816_/A _12601_/B vssd1 vssd1 vccd1 vccd1 _11734_/A sky130_fd_sc_hd__nor2_4
XFILLER_59_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09747_ _18597_/Q _18168_/Q _09770_/S vssd1 vssd1 vccd1 vccd1 _09747_/X sky130_fd_sc_hd__mux2_1
XFILLER_274_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09678_ _10315_/S _09677_/X _10260_/B1 vssd1 vssd1 vccd1 vccd1 _09678_/X sky130_fd_sc_hd__o21a_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ _11640_/A _12647_/B vssd1 vssd1 vccd1 vccd1 _13761_/A sky130_fd_sc_hd__xnor2_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ _11568_/X _11570_/X _11564_/X vssd1 vssd1 vccd1 vccd1 _11571_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_168_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19075_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_183_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13310_ _13330_/B _13312_/A vssd1 vssd1 vccd1 vccd1 _13310_/X sky130_fd_sc_hd__or2_1
XFILLER_195_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10522_ _11279_/B1 _10505_/X _10520_/X _10521_/Y vssd1 vssd1 vccd1 vccd1 _10522_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_14290_ _16608_/A0 _18149_/Q _14301_/S vssd1 vssd1 vccd1 vccd1 _18149_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13241_ _19242_/Q _13425_/A2 _13425_/B1 _19274_/Q vssd1 vssd1 vccd1 vccd1 _13241_/X
+ sky130_fd_sc_hd__a22o_2
X_10453_ _10453_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _10454_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10384_ _10382_/X _10383_/X _08946_/B vssd1 vssd1 vccd1 vccd1 _10384_/X sky130_fd_sc_hd__a21o_1
XFILLER_164_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13172_ _19336_/Q _13246_/A2 _13246_/B1 _19464_/Q _12570_/C vssd1 vssd1 vccd1 vccd1
+ _13172_/X sky130_fd_sc_hd__a221o_1
XFILLER_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ _12219_/A _12128_/C vssd1 vssd1 vccd1 vccd1 _12123_/Y sky130_fd_sc_hd__nor2_1
XFILLER_184_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17980_ _17982_/CLK _17980_/D vssd1 vssd1 vccd1 vccd1 _17980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16931_ _19317_/Q _17184_/B _16947_/S vssd1 vssd1 vccd1 vccd1 _16932_/B sky130_fd_sc_hd__mux2_1
X_12054_ _17902_/Q _12035_/B _12053_/X _12350_/C1 vssd1 vssd1 vccd1 vccd1 _17804_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1800 _17803_/Q vssd1 vssd1 vccd1 vccd1 _12051_/A sky130_fd_sc_hd__buf_4
Xfanout1811 _15718_/C1 vssd1 vssd1 vccd1 vccd1 _14450_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1822 _14340_/A vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__buf_2
XFILLER_104_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1833 fanout1870/X vssd1 vssd1 vccd1 vccd1 _17336_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11005_ _19636_/Q _18925_/Q _11477_/S vssd1 vssd1 vccd1 vccd1 _11005_/X sky130_fd_sc_hd__mux2_1
Xfanout1844 _17322_/A vssd1 vssd1 vccd1 vccd1 _17328_/A sky130_fd_sc_hd__buf_4
XFILLER_237_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16862_ _19300_/Q _17567_/A _16971_/S vssd1 vssd1 vccd1 vccd1 _16863_/B sky130_fd_sc_hd__mux2_1
Xfanout1855 fanout1870/X vssd1 vssd1 vccd1 vccd1 _13987_/C1 sky130_fd_sc_hd__buf_6
X_19650_ _19650_/CLK _19650_/D vssd1 vssd1 vccd1 vccd1 _19650_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1866 _16764_/B1 vssd1 vssd1 vccd1 vccd1 _15946_/C1 sky130_fd_sc_hd__buf_4
XFILLER_277_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1877 _14423_/B vssd1 vssd1 vccd1 vccd1 _17141_/A sky130_fd_sc_hd__buf_6
XFILLER_19_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15813_ _18605_/Q _17703_/A0 _15832_/S vssd1 vssd1 vccd1 vccd1 _18605_/D sky130_fd_sc_hd__mux2_1
Xfanout1888 _16110_/B1 vssd1 vssd1 vccd1 vccd1 _16142_/B1 sky130_fd_sc_hd__buf_4
X_18601_ _18880_/CLK _18601_/D vssd1 vssd1 vccd1 vccd1 _18601_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout890 _13134_/S vssd1 vssd1 vccd1 vccd1 _13130_/A sky130_fd_sc_hd__buf_4
XFILLER_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19581_ _19613_/CLK _19581_/D vssd1 vssd1 vccd1 vccd1 _19581_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1899 _16740_/A vssd1 vssd1 vccd1 vccd1 _16768_/A sky130_fd_sc_hd__buf_4
XFILLER_203_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16793_ _19286_/Q _16794_/B vssd1 vssd1 vccd1 vccd1 _16795_/B sky130_fd_sc_hd__nor2_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18532_ _19197_/CLK _18532_/D vssd1 vssd1 vccd1 vccd1 _18532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15744_ _15744_/A _15744_/B vssd1 vssd1 vccd1 vccd1 _15749_/A sky130_fd_sc_hd__xnor2_2
XFILLER_234_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12956_ _12956_/A _13349_/B vssd1 vssd1 vccd1 vccd1 _12956_/X sky130_fd_sc_hd__and2_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _19642_/CLK _18463_/D vssd1 vssd1 vccd1 vccd1 _18463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11907_ _11833_/Y _11875_/A _11869_/Y _11901_/B _11906_/X vssd1 vssd1 vccd1 vccd1
+ _11908_/B sky130_fd_sc_hd__o221a_4
X_15675_ _17199_/A _15661_/X _15667_/X _15674_/X _15782_/B1 vssd1 vssd1 vccd1 vccd1
+ _15675_/X sky130_fd_sc_hd__a311o_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_250 _18513_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ _12885_/A _13089_/B _13089_/A vssd1 vssd1 vccd1 vccd1 _12888_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_261 input218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_272 input235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _19494_/Q _17423_/B _17412_/X _17413_/Y _17419_/C1 vssd1 vssd1 vccd1 vccd1
+ _19494_/D sky130_fd_sc_hd__o221a_1
X_14626_ _16486_/A0 _18433_/Q _14628_/S vssd1 vssd1 vccd1 vccd1 _18433_/D sky130_fd_sc_hd__mux2_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_283 input246/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11838_ _11859_/B _11783_/Y _11804_/X _14141_/B vssd1 vssd1 vccd1 vccd1 _11838_/X
+ sky130_fd_sc_hd__a22o_1
X_18394_ _19399_/CLK _18394_/D vssd1 vssd1 vccd1 vccd1 _18394_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_260_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_294 _11984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17345_ _19470_/Q _17587_/A _17345_/S vssd1 vssd1 vccd1 vccd1 _17346_/B sky130_fd_sc_hd__mux2_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _18387_/Q _14589_/A2 _14589_/B1 input15/X vssd1 vssd1 vccd1 vccd1 _14558_/B
+ sky130_fd_sc_hd__o22a_1
X_11769_ _18587_/Q _11726_/B _11769_/B1 _11641_/Y vssd1 vssd1 vccd1 vccd1 _11769_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_202_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13508_ _13507_/B _13506_/X _13507_/Y _13930_/B1 _13931_/A vssd1 vssd1 vccd1 vccd1
+ _13508_/X sky130_fd_sc_hd__a221o_1
XFILLER_159_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17276_ _17274_/Y _17275_/X _16048_/A vssd1 vssd1 vccd1 vccd1 _19442_/D sky130_fd_sc_hd__a21oi_1
XFILLER_201_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14488_ _16392_/B _14488_/B _14488_/C vssd1 vssd1 vccd1 vccd1 _17691_/B sky130_fd_sc_hd__and3_4
X_19015_ _19047_/CLK _19015_/D vssd1 vssd1 vccd1 vccd1 _19015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_0__f_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19652_/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16227_ _16426_/A _16260_/B vssd1 vssd1 vccd1 vccd1 _16227_/Y sky130_fd_sc_hd__nand2_1
X_13439_ _13438_/B _13437_/X _13438_/Y _13930_/B1 _13289_/A vssd1 vssd1 vccd1 vccd1
+ _13439_/X sky130_fd_sc_hd__a221o_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16158_ _19425_/Q _15140_/B _14430_/B vssd1 vssd1 vccd1 vccd1 _16158_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15109_ _10061_/X _12318_/A _15426_/B _10027_/A vssd1 vssd1 vccd1 vccd1 _15109_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_115_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08980_ _11513_/A1 _19629_/Q _18918_/Q _11503_/S0 vssd1 vssd1 vccd1 vccd1 _08980_/X
+ sky130_fd_sc_hd__a22o_1
X_16089_ _18747_/Q _16093_/B vssd1 vssd1 vccd1 vccd1 _16089_/Y sky130_fd_sc_hd__nand2_1
XFILLER_130_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09601_ _10371_/S _09600_/X _09599_/X _11199_/S1 vssd1 vssd1 vccd1 vccd1 _09601_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_272_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09532_ _11172_/A1 _18210_/Q _11160_/S _18945_/Q vssd1 vssd1 vccd1 vccd1 _09532_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_237_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ _09461_/X _09462_/X _09463_/S vssd1 vssd1 vccd1 vccd1 _09463_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09394_ _10346_/S _09392_/X _09393_/X _10356_/C1 vssd1 vssd1 vccd1 vccd1 _09394_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_240_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput460 _18120_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[19] sky130_fd_sc_hd__buf_4
XFILLER_267_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput471 _18130_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[29] sky130_fd_sc_hd__buf_4
XFILLER_248_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput482 _12461_/A vssd1 vssd1 vccd1 vccd1 probe_state sky130_fd_sc_hd__buf_4
XFILLER_78_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_182_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17951_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout1107 _12588_/Y vssd1 vssd1 vccd1 vccd1 _13253_/B1 sky130_fd_sc_hd__buf_2
Xfanout1118 _13968_/B2 vssd1 vssd1 vccd1 vccd1 _13323_/B sky130_fd_sc_hd__buf_4
XFILLER_232_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1129 _12323_/X vssd1 vssd1 vccd1 vccd1 _15124_/B sky130_fd_sc_hd__buf_4
XFILLER_232_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_111_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19276_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_247_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12810_ _12810_/A vssd1 vssd1 vccd1 vccd1 _12810_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13790_ _13758_/A _13775_/X _13956_/B1 vssd1 vssd1 vccd1 vccd1 _13791_/C sky130_fd_sc_hd__a21o_1
XFILLER_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12445_/B _12740_/X _09075_/X vssd1 vssd1 vccd1 vccd1 _12741_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15460_ _15407_/X _15430_/Y _15431_/Y _15459_/X vssd1 vssd1 vccd1 vccd1 _15460_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_179_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12672_ _09401_/C _12729_/B _12671_/X vssd1 vssd1 vccd1 vccd1 _12672_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_179_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14411_ _17718_/A0 _18262_/Q _14416_/S vssd1 vssd1 vccd1 vccd1 _18262_/D sky130_fd_sc_hd__mux2_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11623_/A1 _11621_/X _11622_/X _11608_/X vssd1 vssd1 vccd1 vccd1 _11623_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_230_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15391_ _15391_/A _15456_/B vssd1 vssd1 vccd1 vccd1 _15391_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_169_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17130_ _08881_/X _15118_/B _17129_/Y vssd1 vssd1 vccd1 vccd1 _17130_/Y sky130_fd_sc_hd__a21oi_1
X_14342_ _14342_/A _14345_/B _14342_/C vssd1 vssd1 vccd1 vccd1 _18197_/D sky130_fd_sc_hd__and3_4
XFILLER_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11554_ _10232_/Y _11636_/A _11553_/B _11634_/B vssd1 vssd1 vccd1 vccd1 _11555_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17061_ _19364_/Q _17073_/B vssd1 vssd1 vccd1 vccd1 _17061_/X sky130_fd_sc_hd__or2_1
X_10505_ _11131_/A _10499_/X _10502_/X _10504_/X vssd1 vssd1 vccd1 vccd1 _10505_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14273_ _16260_/B _17691_/A vssd1 vssd1 vccd1 vccd1 _14273_/Y sky130_fd_sc_hd__nand2_2
X_11485_ _11463_/X _11466_/X _11484_/X vssd1 vssd1 vccd1 vccd1 _11485_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_155_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _18721_/Q _15953_/B _16147_/A2 _18770_/Q _16018_/C1 vssd1 vssd1 vccd1 vccd1
+ _16012_/X sky130_fd_sc_hd__a221o_1
X_13224_ _13224_/A _13224_/B vssd1 vssd1 vccd1 vccd1 _13224_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10436_ _10434_/X _10435_/X _11606_/S vssd1 vssd1 vccd1 vccd1 _10436_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13155_ _14156_/A0 _13154_/X _09403_/B vssd1 vssd1 vccd1 vccd1 _13155_/Y sky130_fd_sc_hd__o21ai_4
X_10367_ _10364_/X _10365_/X _10366_/X _10742_/A1 _10746_/S vssd1 vssd1 vccd1 vccd1
+ _10367_/X sky130_fd_sc_hd__a221o_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _17828_/Q _17829_/Q _12106_/C vssd1 vssd1 vccd1 vccd1 _12112_/C sky130_fd_sc_hd__and3_2
XFILLER_152_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17963_ _17982_/CLK _17963_/D vssd1 vssd1 vccd1 vccd1 _17963_/Q sky130_fd_sc_hd__dfxtp_1
X_10298_ _18467_/Q _18368_/Q _10299_/S vssd1 vssd1 vccd1 vccd1 _10298_/X sky130_fd_sc_hd__mux2_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _12874_/X _12885_/Y _13089_/A vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1630 _12024_/A vssd1 vssd1 vccd1 vccd1 _09062_/B sky130_fd_sc_hd__buf_6
X_16914_ _16848_/S _17937_/Q _16913_/X vssd1 vssd1 vccd1 vccd1 _17172_/B sky130_fd_sc_hd__o21a_4
X_12037_ _17796_/Q _12051_/B vssd1 vssd1 vccd1 vccd1 _12037_/X sky130_fd_sc_hd__or2_1
XFILLER_66_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1641 _11596_/A1 vssd1 vssd1 vccd1 vccd1 _11360_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_266_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17894_ _17958_/CLK _17894_/D vssd1 vssd1 vccd1 vccd1 _17894_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1652 _10282_/A1 vssd1 vssd1 vccd1 vccd1 _10366_/A1 sky130_fd_sc_hd__buf_6
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1663 _10030_/C1 vssd1 vssd1 vccd1 vccd1 _08899_/A sky130_fd_sc_hd__buf_12
Xfanout1674 _08846_/Y vssd1 vssd1 vccd1 vccd1 _11607_/S sky130_fd_sc_hd__buf_12
Xfanout1685 _08845_/Y vssd1 vssd1 vccd1 vccd1 _10625_/A1 sky130_fd_sc_hd__buf_8
X_19633_ _19640_/CLK _19633_/D vssd1 vssd1 vccd1 vccd1 _19633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16845_ _16846_/B vssd1 vssd1 vccd1 vccd1 _17117_/B sky130_fd_sc_hd__inv_2
XFILLER_93_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1696 _11458_/A1 vssd1 vssd1 vccd1 vccd1 _11465_/A1 sky130_fd_sc_hd__buf_4
XFILLER_225_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19564_ _19564_/CLK _19564_/D vssd1 vssd1 vccd1 vccd1 _19564_/Q sky130_fd_sc_hd__dfxtp_1
X_16776_ _16776_/A _16776_/B _16778_/B vssd1 vssd1 vccd1 vccd1 _19279_/D sky130_fd_sc_hd__nor3_1
XFILLER_280_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13988_ _14020_/B _13988_/B vssd1 vssd1 vccd1 vccd1 _13988_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18515_ _18517_/CLK _18515_/D vssd1 vssd1 vccd1 vccd1 _18515_/Q sky130_fd_sc_hd__dfxtp_4
X_15727_ _15644_/B _15685_/A _15686_/X _15707_/A _15726_/Y vssd1 vssd1 vccd1 vccd1
+ _15728_/B sky130_fd_sc_hd__o41a_2
XFILLER_280_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12939_ _12942_/S _12804_/X _12938_/Y vssd1 vssd1 vccd1 vccd1 _13129_/B sky130_fd_sc_hd__o21ai_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19495_ _19526_/CLK _19495_/D vssd1 vssd1 vccd1 vccd1 _19495_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18446_ _19625_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_1
X_15658_ _18126_/Q _15763_/A2 _15657_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _15687_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14609_ _16535_/A0 _18416_/Q _14630_/S vssd1 vssd1 vccd1 vccd1 _18416_/D sky130_fd_sc_hd__mux2_1
X_18377_ _19471_/CLK _18377_/D vssd1 vssd1 vccd1 vccd1 _18377_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15589_ _19477_/Q _19411_/Q vssd1 vssd1 vccd1 vccd1 _15590_/B sky130_fd_sc_hd__nor2_1
XFILLER_175_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17328_ _17328_/A _17328_/B vssd1 vssd1 vccd1 vccd1 _19461_/D sky130_fd_sc_hd__and2_1
XFILLER_239_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17259_ _17457_/A _17250_/B _18114_/Q _17129_/A vssd1 vssd1 vccd1 vccd1 _17259_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_174_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08963_ _10427_/C1 _08962_/X _11417_/B1 vssd1 vssd1 vccd1 vccd1 _08963_/X sky130_fd_sc_hd__a21o_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08894_ _10373_/S _09285_/C vssd1 vssd1 vccd1 vccd1 _08894_/Y sky130_fd_sc_hd__nand2_8
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09515_ _19105_/Q _19137_/Q _09883_/B vssd1 vssd1 vccd1 vccd1 _09515_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09446_ _18414_/Q _11167_/B _09445_/X _10264_/S vssd1 vssd1 vccd1 vccd1 _09446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09377_ _10373_/S _09374_/X _09376_/Y _09958_/C1 vssd1 vssd1 vccd1 vccd1 _09377_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_197_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11270_ _11268_/X _11269_/X _11285_/S vssd1 vssd1 vccd1 vccd1 _11270_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10221_ _09708_/A _10216_/X _10220_/X _08895_/A vssd1 vssd1 vccd1 vccd1 _10221_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10152_ _10148_/X _10151_/X _10301_/S vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput290 _11965_/X vssd1 vssd1 vccd1 vccd1 addr0[5] sky130_fd_sc_hd__buf_4
X_10083_ _11556_/C _09025_/A _09025_/B _09987_/A vssd1 vssd1 vccd1 vccd1 _10083_/X
+ sky130_fd_sc_hd__a31o_1
X_14960_ _14956_/Y _14959_/X _15010_/B1 vssd1 vssd1 vccd1 vccd1 _14960_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13911_ _13911_/A _13911_/B vssd1 vssd1 vccd1 vccd1 _13911_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14891_ _15003_/A1 _13594_/Y _15003_/B1 _18646_/Q _15003_/C1 vssd1 vssd1 vccd1 vccd1
+ _14891_/X sky130_fd_sc_hd__a221o_1
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16630_ _17724_/A _19232_/Q _16752_/A vssd1 vssd1 vccd1 vccd1 _16630_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13842_ _17947_/Q _13940_/A2 _13841_/X _14181_/A vssd1 vssd1 vccd1 vccd1 _17947_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16561_ _16594_/A0 _19165_/Q _16586_/S vssd1 vssd1 vccd1 vccd1 _19165_/D sky130_fd_sc_hd__mux2_1
XFILLER_244_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13773_ _17913_/Q _12448_/C _12762_/B _13772_/Y vssd1 vssd1 vccd1 vccd1 _13773_/X
+ sky130_fd_sc_hd__a211o_4
X_10985_ _10985_/A _10985_/B vssd1 vssd1 vccd1 vccd1 _11673_/B sky130_fd_sc_hd__or2_4
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18300_ _19450_/CLK _18300_/D vssd1 vssd1 vccd1 vccd1 _18300_/Q sky130_fd_sc_hd__dfxtp_1
X_15512_ _18580_/Q _18579_/Q _15512_/C vssd1 vssd1 vccd1 vccd1 _15561_/C sky130_fd_sc_hd__and3_2
XFILLER_71_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19280_ _19280_/CLK _19280_/D vssd1 vssd1 vccd1 vccd1 _19280_/Q sky130_fd_sc_hd__dfxtp_1
X_12724_ _11136_/Y _12596_/B _12729_/B vssd1 vssd1 vccd1 vccd1 _12823_/B sky130_fd_sc_hd__mux2_1
X_16492_ _16525_/A _17691_/A vssd1 vssd1 vccd1 vccd1 _16492_/Y sky130_fd_sc_hd__nand2_8
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18231_ _19596_/CLK _18231_/D vssd1 vssd1 vccd1 vccd1 _18231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15443_ _19471_/Q _19405_/Q vssd1 vssd1 vccd1 vccd1 _15444_/B sky130_fd_sc_hd__or2_1
X_12655_ _11639_/A _13727_/B _12647_/Y _12654_/Y vssd1 vssd1 vccd1 vccd1 _13860_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_230_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18162_ _19193_/CLK _18162_/D vssd1 vssd1 vccd1 vccd1 _18162_/Q sky130_fd_sc_hd__dfxtp_1
X_11606_ _11604_/X _11605_/X _11606_/S vssd1 vssd1 vccd1 vccd1 _11606_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15374_ _19467_/Q _19401_/Q _15347_/B vssd1 vssd1 vccd1 vccd1 _15374_/X sky130_fd_sc_hd__a21o_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12586_ _12756_/B _12587_/B vssd1 vssd1 vccd1 vccd1 _12586_/X sky130_fd_sc_hd__and2_4
XFILLER_184_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17113_ _19390_/Q _17113_/B vssd1 vssd1 vccd1 vccd1 _17113_/X sky130_fd_sc_hd__or2_1
X_14325_ _18182_/Q _17676_/A0 _14325_/S vssd1 vssd1 vccd1 vccd1 _18182_/D sky130_fd_sc_hd__mux2_1
X_18093_ _19306_/CLK _18093_/D vssd1 vssd1 vccd1 vccd1 _18093_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11537_ _11537_/A _11537_/B vssd1 vssd1 vccd1 vccd1 _13616_/A sky130_fd_sc_hd__nor2_8
XFILLER_129_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17044_ _17211_/B _17044_/A2 _17043_/X _17378_/A vssd1 vssd1 vccd1 vccd1 _19358_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14256_ _18126_/Q _14260_/B vssd1 vssd1 vccd1 vccd1 _14256_/X sky130_fd_sc_hd__or2_1
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11468_ _18352_/Q _10101_/B _11467_/X vssd1 vssd1 vccd1 vccd1 _11468_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_171_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13207_ _19241_/Q _13425_/A2 _13425_/B1 _19273_/Q vssd1 vssd1 vccd1 vccd1 _13207_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10419_ _10417_/X _10418_/X _10419_/S vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__mux2_1
X_14187_ _16972_/A _14187_/B vssd1 vssd1 vccd1 vccd1 _18091_/D sky130_fd_sc_hd__and2_1
X_11399_ _18824_/Q _11479_/B vssd1 vssd1 vccd1 vccd1 _11399_/X sky130_fd_sc_hd__or2_1
XFILLER_125_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13138_ _13414_/A _12719_/B _12745_/X vssd1 vssd1 vccd1 vccd1 _13139_/A sky130_fd_sc_hd__o21a_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _19611_/CLK _18995_/D vssd1 vssd1 vccd1 vccd1 _18995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _18627_/CLK _17946_/D vssd1 vssd1 vccd1 vccd1 _17946_/Q sky130_fd_sc_hd__dfxtp_2
X_13069_ _13246_/B1 _13243_/B1 _12570_/X _12568_/Y _19489_/Q vssd1 vssd1 vccd1 vccd1
+ _13069_/X sky130_fd_sc_hd__o32a_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1460 _10217_/B vssd1 vssd1 vccd1 vccd1 _10364_/B sky130_fd_sc_hd__buf_12
XFILLER_39_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1471 _10656_/S vssd1 vssd1 vccd1 vccd1 _10582_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17877_ _19319_/CLK _17877_/D vssd1 vssd1 vccd1 vccd1 _17877_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1482 fanout1485/X vssd1 vssd1 vccd1 vccd1 _10744_/S sky130_fd_sc_hd__clkbuf_8
Xfanout1493 _10721_/S vssd1 vssd1 vccd1 vccd1 _09720_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_253_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19616_ _19648_/CLK _19616_/D vssd1 vssd1 vccd1 vccd1 _19616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16828_ _16973_/B _17118_/B vssd1 vssd1 vccd1 vccd1 _17217_/A sky130_fd_sc_hd__nand2b_1
XFILLER_254_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19547_ _19553_/CLK _19547_/D vssd1 vssd1 vccd1 vccd1 _19547_/Q sky130_fd_sc_hd__dfxtp_1
X_16759_ _19273_/Q _19272_/Q _16759_/C vssd1 vssd1 vccd1 vccd1 _16762_/B sky130_fd_sc_hd__and3_1
XFILLER_0_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09300_ _09298_/X _09299_/X _09967_/S vssd1 vssd1 vccd1 vccd1 _09300_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19478_ _19483_/CLK _19478_/D vssd1 vssd1 vccd1 vccd1 _19478_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09231_ input124/X input159/X _09655_/S vssd1 vssd1 vccd1 vccd1 _09232_/B sky130_fd_sc_hd__mux2_8
XFILLER_221_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18429_ _19146_/CLK _18429_/D vssd1 vssd1 vccd1 vccd1 _18429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09162_ _18853_/Q _18885_/Q _10099_/S vssd1 vssd1 vccd1 vccd1 _09162_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09093_ _09457_/B _09285_/C vssd1 vssd1 vccd1 vccd1 _09093_/Y sky130_fd_sc_hd__nand2_4
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09995_ _08946_/B _09988_/Y _09994_/X _17920_/Q vssd1 vssd1 vccd1 vccd1 _09995_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_130_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08946_ _08947_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _08946_/Y sky130_fd_sc_hd__nor2_8
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08877_ _17917_/Q _17916_/Q _17915_/Q vssd1 vssd1 vccd1 vccd1 _09073_/D sky130_fd_sc_hd__or3_4
XFILLER_229_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10770_ _10768_/X _10769_/X _11577_/S vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ _09427_/X _09428_/X _09429_/S vssd1 vssd1 vccd1 vccd1 _09429_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12440_ _12756_/A _12455_/A vssd1 vssd1 vccd1 vccd1 _12440_/X sky130_fd_sc_hd__and2_2
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12371_ _17898_/Q _12382_/A _12370_/Y _12383_/C1 vssd1 vssd1 vccd1 vccd1 _17898_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14110_ _16461_/A0 _18049_/Q _14137_/S vssd1 vssd1 vccd1 vccd1 _18049_/D sky130_fd_sc_hd__mux2_1
X_11322_ _18250_/Q _18825_/Q _11325_/S vssd1 vssd1 vccd1 vccd1 _11322_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15090_ _19385_/Q _15092_/B _15090_/C vssd1 vssd1 vccd1 vccd1 _15093_/C sky130_fd_sc_hd__and3_1
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14041_ _17658_/A _16393_/A vssd1 vssd1 vccd1 vccd1 _14041_/Y sky130_fd_sc_hd__nand2_8
XFILLER_107_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11253_ _11227_/X _11230_/X _10326_/A vssd1 vssd1 vccd1 vccd1 _11253_/X sky130_fd_sc_hd__a21o_1
XFILLER_180_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10204_ _19128_/Q _19160_/Q _10206_/S vssd1 vssd1 vccd1 vccd1 _10204_/X sky130_fd_sc_hd__mux2_1
X_11184_ _08901_/A _19634_/Q _18923_/Q _09883_/B vssd1 vssd1 vccd1 vccd1 _11184_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17800_ _18201_/CLK _17800_/D vssd1 vssd1 vccd1 vccd1 _17800_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_122_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10135_ _10200_/S _10127_/X _10126_/X _10356_/C1 vssd1 vssd1 vccd1 vccd1 _10135_/X
+ sky130_fd_sc_hd__a211o_1
X_15992_ _18711_/Q _16002_/A2 _16004_/B1 _18760_/Q _16004_/C1 vssd1 vssd1 vccd1 vccd1
+ _15992_/X sky130_fd_sc_hd__a221o_1
X_18780_ _19619_/CLK _18780_/D vssd1 vssd1 vccd1 vccd1 _18780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17731_ _18631_/Q vssd1 vssd1 vccd1 vccd1 _18631_/D sky130_fd_sc_hd__clkbuf_2
X_10066_ _12838_/S _11653_/A vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__nor2_4
X_14943_ _15003_/A1 _13756_/Y _15003_/B1 _18651_/Q _15003_/C1 vssd1 vssd1 vccd1 vccd1
+ _14943_/X sky130_fd_sc_hd__a221o_1
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14874_ _18119_/Q _14801_/B _14852_/X _14873_/X vssd1 vssd1 vccd1 vccd1 _14874_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17662_ _17662_/A0 _19589_/Q _17681_/S vssd1 vssd1 vccd1 vccd1 _19589_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19401_ _19433_/CLK _19401_/D vssd1 vssd1 vccd1 vccd1 _19401_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_263_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16613_ _17713_/A0 _19216_/Q _16618_/S vssd1 vssd1 vccd1 vccd1 _19216_/D sky130_fd_sc_hd__mux2_1
X_13825_ _19419_/Q _13948_/A2 _13948_/B1 vssd1 vssd1 vccd1 vccd1 _13825_/X sky130_fd_sc_hd__a21o_1
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17593_ _19376_/Q _15086_/B input171/X _17592_/X _17623_/B1 vssd1 vssd1 vccd1 vccd1
+ _17593_/X sky130_fd_sc_hd__a41o_1
XFILLER_251_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16544_ _17644_/A0 _19149_/Q _16556_/S vssd1 vssd1 vccd1 vccd1 _19149_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19332_ _19526_/CLK _19332_/D vssd1 vssd1 vccd1 vccd1 _19332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13756_ _14024_/B vssd1 vssd1 vccd1 vccd1 _13756_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10968_ _11358_/A _10967_/X _11608_/C1 vssd1 vssd1 vccd1 vccd1 _10968_/X sky130_fd_sc_hd__a21o_1
X_12707_ _12603_/B _13911_/A _12743_/A vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__a21bo_1
X_19263_ _19295_/CLK _19263_/D vssd1 vssd1 vccd1 vccd1 _19263_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16475_ _17674_/A0 _19082_/Q _16485_/S vssd1 vssd1 vccd1 vccd1 _19082_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13687_ _19447_/Q _13949_/A2 _13685_/X _13686_/X _13949_/C1 vssd1 vssd1 vccd1 vccd1
+ _13687_/X sky130_fd_sc_hd__o221a_1
XFILLER_188_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10899_ _11112_/A _10894_/X _10898_/X vssd1 vssd1 vccd1 vccd1 _10901_/C sky130_fd_sc_hd__a21oi_1
XFILLER_15_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18214_ _19564_/CLK _18214_/D vssd1 vssd1 vccd1 vccd1 _18214_/Q sky130_fd_sc_hd__dfxtp_1
X_15426_ _15426_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15426_/X sky130_fd_sc_hd__and2_1
X_12638_ _12638_/A _13597_/A _13616_/A _13697_/A vssd1 vssd1 vccd1 vccd1 _12638_/Y
+ sky130_fd_sc_hd__nor4_1
X_19194_ _19226_/CLK _19194_/D vssd1 vssd1 vccd1 vccd1 _19194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18145_ _19208_/CLK _18145_/D vssd1 vssd1 vccd1 vccd1 _18145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15357_ _15357_/A _15404_/B vssd1 vssd1 vccd1 vccd1 _15357_/Y sky130_fd_sc_hd__nor2_1
XFILLER_184_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12569_ _12552_/A _12580_/A _12562_/B vssd1 vssd1 vccd1 vccd1 _12569_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14308_ _18165_/Q _16592_/A0 _14325_/S vssd1 vssd1 vccd1 vccd1 _18165_/D sky130_fd_sc_hd__mux2_1
X_18076_ _19626_/CLK _18076_/D vssd1 vssd1 vccd1 vccd1 _18076_/Q sky130_fd_sc_hd__dfxtp_1
X_15288_ _15289_/A _15289_/B vssd1 vssd1 vccd1 vccd1 _15290_/A sky130_fd_sc_hd__nand2_1
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17027_ _19350_/Q _17045_/B vssd1 vssd1 vccd1 vccd1 _17027_/X sky130_fd_sc_hd__or2_1
X_14239_ _18291_/Q _14267_/A2 _14238_/X _14452_/B vssd1 vssd1 vccd1 vccd1 _18117_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout708 _12543_/X vssd1 vssd1 vccd1 vccd1 _13105_/B sky130_fd_sc_hd__buf_2
XFILLER_259_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout719 _12532_/Y vssd1 vssd1 vccd1 vccd1 _13952_/A2 sky130_fd_sc_hd__buf_8
XFILLER_213_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09780_ _18104_/Q _09948_/B vssd1 vssd1 vccd1 vccd1 _09780_/X sky130_fd_sc_hd__or2_1
X_18978_ _19138_/CLK _18978_/D vssd1 vssd1 vccd1 vccd1 _18978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17929_ _17931_/CLK _17929_/D vssd1 vssd1 vccd1 vccd1 _17929_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1290 _15014_/Y vssd1 vssd1 vccd1 vccd1 _15037_/S sky130_fd_sc_hd__buf_6
XFILLER_227_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ _18026_/Q _17994_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _09214_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09145_ _09145_/A _13267_/A vssd1 vssd1 vccd1 vccd1 _13261_/A sky130_fd_sc_hd__nor2_4
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09076_ _12442_/A _12837_/A _12443_/B vssd1 vssd1 vccd1 vccd1 _12740_/C sky130_fd_sc_hd__a21o_1
XFILLER_190_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18700_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09978_ _09978_/A1 _09972_/X _09975_/X _08904_/A vssd1 vssd1 vccd1 vccd1 _09978_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19114_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08929_ _08940_/B _08929_/B _08942_/B _08929_/D vssd1 vssd1 vccd1 vccd1 _08929_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_258_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _11944_/A1 _11857_/B _11945_/B1 input227/X vssd1 vssd1 vccd1 vccd1 _11940_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_206_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11871_ _14141_/B _11833_/Y _11869_/Y _11952_/A2 _11870_/X vssd1 vssd1 vccd1 vccd1
+ _11872_/B sky130_fd_sc_hd__a221oi_4
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _13904_/A _13610_/B vssd1 vssd1 vccd1 vccd1 _13610_/Y sky130_fd_sc_hd__nand2_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _10820_/X _10821_/X _11606_/S vssd1 vssd1 vccd1 vccd1 _10822_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14592_/A _14590_/B vssd1 vssd1 vccd1 vccd1 _18403_/D sky130_fd_sc_hd__or2_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13541_ _18119_/Q _13541_/B vssd1 vssd1 vccd1 vccd1 _13542_/B sky130_fd_sc_hd__nor2_1
XFILLER_241_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10753_ _10753_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _10754_/B sky130_fd_sc_hd__nor2_4
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16260_ _16393_/A _16260_/B vssd1 vssd1 vccd1 vccd1 _16260_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13472_ _12447_/Y _13471_/X _13463_/X vssd1 vssd1 vccd1 vccd1 _13472_/X sky130_fd_sc_hd__a21bo_1
XFILLER_201_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ _19640_/Q _18929_/Q _11249_/S vssd1 vssd1 vccd1 vccd1 _10684_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15211_ _17382_/A _15205_/X _15210_/X _15424_/C1 vssd1 vssd1 vccd1 vccd1 _15211_/X
+ sky130_fd_sc_hd__a211o_1
X_12423_ _12429_/A1 _09232_/A _09655_/X _12429_/B1 _18401_/Q vssd1 vssd1 vccd1 vccd1
+ _12424_/B sky130_fd_sc_hd__o32ai_4
X_16191_ _16621_/A0 _18808_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _18808_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15142_ _19392_/Q _15400_/S _19458_/Q vssd1 vssd1 vccd1 vccd1 _15145_/B sky130_fd_sc_hd__a21oi_1
X_12354_ _11695_/B _09991_/A _09563_/X _12432_/B1 _18378_/Q vssd1 vssd1 vccd1 vccd1
+ _12355_/B sky130_fd_sc_hd__o32ai_2
XFILLER_193_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11305_ _11305_/A1 _19145_/Q _11302_/S _19113_/Q _10784_/S vssd1 vssd1 vccd1 vccd1
+ _11305_/X sky130_fd_sc_hd__o221a_1
X_15073_ _18557_/Q _16551_/A0 _15079_/S vssd1 vssd1 vccd1 vccd1 _18557_/D sky130_fd_sc_hd__mux2_1
X_12285_ _12285_/A _12478_/B _12492_/B _12284_/X vssd1 vssd1 vccd1 vccd1 _14688_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14024_ _14028_/A _14024_/B vssd1 vssd1 vccd1 vccd1 _14024_/Y sky130_fd_sc_hd__nand2_1
X_18901_ _19055_/CLK _18901_/D vssd1 vssd1 vccd1 vccd1 _18901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11236_ _11565_/A1 _17773_/Q _11247_/S _18322_/Q _11567_/S vssd1 vssd1 vccd1 vccd1
+ _11236_/X sky130_fd_sc_hd__o221a_1
XFILLER_267_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18832_ _19639_/CLK _18832_/D vssd1 vssd1 vccd1 vccd1 _18832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11167_ _18827_/Q _11167_/B vssd1 vssd1 vccd1 vccd1 _11167_/X sky130_fd_sc_hd__or2_1
XFILLER_110_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10118_ _10115_/X _10117_/X _11484_/B1 vssd1 vssd1 vccd1 vccd1 _10118_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18763_ _18772_/CLK _18763_/D vssd1 vssd1 vccd1 vccd1 _18763_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_212_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ _18703_/Q _16003_/A2 _15974_/X _16972_/A vssd1 vssd1 vccd1 vccd1 _18703_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_209_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11098_ _11071_/X _11074_/X _10399_/A vssd1 vssd1 vccd1 vccd1 _11098_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17714_ _17714_/A0 _19640_/Q _17719_/S vssd1 vssd1 vccd1 vccd1 _19640_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14926_ input58/X input93/X _14947_/S vssd1 vssd1 vccd1 vccd1 _14927_/A sky130_fd_sc_hd__mux2_2
X_10049_ _18016_/Q _17984_/Q _10726_/S vssd1 vssd1 vccd1 vccd1 _10049_/X sky130_fd_sc_hd__mux2_1
X_18694_ _18749_/CLK _18694_/D vssd1 vssd1 vccd1 vccd1 _18694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17645_ _17678_/A0 _19573_/Q _17657_/S vssd1 vssd1 vccd1 vccd1 _19573_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14857_ _14857_/A vssd1 vssd1 vccd1 vccd1 _14857_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13808_ _17914_/Q _12762_/A _13806_/Y _13807_/X _13808_/C1 vssd1 vssd1 vccd1 vccd1
+ _13808_/X sky130_fd_sc_hd__a221o_4
X_14788_ _18480_/Q _14889_/B1 _14787_/Y _12243_/A vssd1 vssd1 vccd1 vccd1 _18480_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17576_ _19530_/Q _17561_/B _17588_/B1 _17575_/X vssd1 vssd1 vccd1 vccd1 _19530_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19315_ _19363_/CLK _19315_/D vssd1 vssd1 vccd1 vccd1 _19315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16527_ _17660_/A0 _19132_/Q _16554_/S vssd1 vssd1 vccd1 vccd1 _19132_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13739_ _13739_/A _13739_/B vssd1 vssd1 vccd1 vccd1 _13739_/Y sky130_fd_sc_hd__nand2_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19246_ _19280_/CLK _19246_/D vssd1 vssd1 vccd1 vccd1 _19246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16458_ _19066_/Q _17723_/A0 _16458_/S vssd1 vssd1 vccd1 vccd1 _19066_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409_ _15385_/A _15385_/B _15386_/Y _15384_/Y vssd1 vssd1 vccd1 vccd1 _15410_/B
+ sky130_fd_sc_hd__a31o_1
X_16389_ _16522_/A0 _19000_/Q _16390_/S vssd1 vssd1 vccd1 vccd1 _19000_/D sky130_fd_sc_hd__mux2_1
XFILLER_191_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19177_ _19632_/CLK _19177_/D vssd1 vssd1 vccd1 vccd1 _19177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18128_ _19450_/CLK _18128_/D vssd1 vssd1 vccd1 vccd1 _18128_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_247_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18059_ _19140_/CLK _18059_/D vssd1 vssd1 vccd1 vccd1 _18059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ _09901_/A _11556_/B _09000_/Y vssd1 vssd1 vccd1 vccd1 _09903_/C sky130_fd_sc_hd__or3b_1
XFILLER_259_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout505 _11706_/X vssd1 vssd1 vccd1 vccd1 _14667_/A1 sky130_fd_sc_hd__buf_8
Xfanout516 _17219_/Y vssd1 vssd1 vccd1 vccd1 _17313_/B sky130_fd_sc_hd__buf_6
XFILLER_99_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout527 _11729_/X vssd1 vssd1 vccd1 vccd1 _11769_/B1 sky130_fd_sc_hd__buf_8
X_09832_ _11157_/A1 _18596_/Q _18167_/Q _10001_/S vssd1 vssd1 vccd1 vccd1 _09832_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_258_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout538 _15499_/B1 vssd1 vssd1 vccd1 vccd1 _15424_/C1 sky130_fd_sc_hd__buf_6
XFILLER_59_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout549 _17199_/A vssd1 vssd1 vccd1 vccd1 _17208_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09763_ _09761_/X _09762_/X _11562_/S vssd1 vssd1 vccd1 vccd1 _09764_/B sky130_fd_sc_hd__mux2_1
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09694_ _09611_/A _09662_/X _09693_/Y vssd1 vssd1 vccd1 vccd1 _11793_/B sky130_fd_sc_hd__o21ai_4
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_136_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19326_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09128_ _18247_/Q _18822_/Q _18450_/Q _18351_/Q _09269_/S _12466_/A0 vssd1 vssd1
+ vccd1 vccd1 _09128_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09059_ _17901_/Q _12442_/B vssd1 vssd1 vccd1 vccd1 _12264_/A sky130_fd_sc_hd__nand2_8
XFILLER_123_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12070_ _15129_/B2 _12088_/A2 _12069_/X _17419_/C1 vssd1 vssd1 vccd1 vccd1 _17812_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11021_ _11000_/X _11003_/X _11020_/X vssd1 vssd1 vccd1 vccd1 _11021_/X sky130_fd_sc_hd__a21o_1
XFILLER_173_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _15751_/X _15752_/X _15759_/X _15782_/A1 _15782_/B1 vssd1 vssd1 vccd1 vccd1
+ _15760_/X sky130_fd_sc_hd__a221o_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _19332_/Q _13246_/A2 _13246_/B1 _19460_/Q _12570_/C vssd1 vssd1 vccd1 vccd1
+ _12972_/X sky130_fd_sc_hd__a221o_1
XFILLER_64_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _18472_/Q _14720_/A _14710_/Y _17330_/A vssd1 vssd1 vccd1 vccd1 _18472_/D
+ sky130_fd_sc_hd__a211o_1
X_11923_ _11926_/A1 _11939_/A1 wire989/X _11935_/B1 input240/X vssd1 vssd1 vccd1 vccd1
+ _11923_/X sky130_fd_sc_hd__a32o_4
XFILLER_245_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _19450_/Q _15793_/A2 _15679_/X _15690_/Y _17199_/A vssd1 vssd1 vccd1 vccd1
+ _15691_/X sky130_fd_sc_hd__o221a_1
XFILLER_73_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_410 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_421 _13810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14642_ _17701_/A0 _18448_/Q _14663_/S vssd1 vssd1 vccd1 vccd1 _18448_/D sky130_fd_sc_hd__mux2_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_432 _11849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _13147_/A _17445_/A2 _17445_/B1 _17798_/Q _17445_/C1 vssd1 vssd1 vccd1 vccd1
+ _17430_/X sky130_fd_sc_hd__a221o_1
XANTENNA_443 _14000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ _11854_/A _11864_/B vssd1 vssd1 vccd1 vccd1 _11854_/X sky130_fd_sc_hd__or2_2
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_454 _19390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_465 _18374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_476 input223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10805_ _11594_/A1 _18225_/Q _11604_/S _18960_/Q _11355_/A1 vssd1 vssd1 vccd1 vccd1
+ _10805_/X sky130_fd_sc_hd__o221a_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_487 _18734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17361_ _19478_/Q _17187_/B _17361_/S vssd1 vssd1 vccd1 vccd1 _17362_/B sky130_fd_sc_hd__mux2_1
X_14573_ _18395_/Q _14575_/A2 _14575_/B1 input24/X vssd1 vssd1 vccd1 vccd1 _14574_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_498 _14277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ _11816_/A _11785_/B vssd1 vssd1 vccd1 vccd1 _11807_/B sky130_fd_sc_hd__nor2_8
X_19100_ _19587_/CLK _19100_/D vssd1 vssd1 vccd1 vccd1 _19100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16312_ _17710_/A0 _18925_/Q _16324_/S vssd1 vssd1 vccd1 vccd1 _18925_/D sky130_fd_sc_hd__mux2_1
X_13524_ _19346_/Q _13883_/A2 _13883_/B1 _19474_/Q _13883_/C1 vssd1 vssd1 vccd1 vccd1
+ _13524_/X sky130_fd_sc_hd__a221o_1
XFILLER_242_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17292_ _19448_/Q _17307_/B vssd1 vssd1 vccd1 vccd1 _17292_/Y sky130_fd_sc_hd__nand2_1
X_10736_ _10732_/X _10733_/X _10745_/S vssd1 vssd1 vccd1 vccd1 _10736_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19031_ _19625_/CLK _19031_/D vssd1 vssd1 vccd1 vccd1 _19031_/Q sky130_fd_sc_hd__dfxtp_1
X_16243_ _16607_/A0 _18858_/Q _16245_/S vssd1 vssd1 vccd1 vccd1 _18858_/D sky130_fd_sc_hd__mux2_1
X_13455_ _19344_/Q _13950_/A2 _13950_/B1 _19472_/Q _13950_/C1 vssd1 vssd1 vccd1 vccd1
+ _13455_/X sky130_fd_sc_hd__a221o_1
X_10667_ _19641_/Q _18930_/Q _10667_/S vssd1 vssd1 vccd1 vccd1 _10667_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12406_ _12430_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _12406_/Y sky130_fd_sc_hd__nand2_1
X_16174_ _11452_/B _18791_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _18791_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13386_ _13351_/A _13351_/B _12597_/Y vssd1 vssd1 vccd1 vccd1 _13387_/B sky130_fd_sc_hd__o21ba_1
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10598_ _11365_/B2 _16418_/A0 _10597_/X _11133_/B2 vssd1 vssd1 vccd1 vccd1 _13711_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_15125_ _17211_/A _15731_/B1 _14224_/B vssd1 vssd1 vccd1 vccd1 _16156_/B sky130_fd_sc_hd__a21o_2
X_12337_ _17887_/Q _14224_/B _12336_/X _14423_/B vssd1 vssd1 vccd1 vccd1 _17887_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15056_ _18540_/Q _16501_/A0 _15078_/S vssd1 vssd1 vccd1 vccd1 _18540_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12268_ _09080_/C _13227_/C1 _12314_/B _12263_/A vssd1 vssd1 vccd1 vccd1 _15082_/C
+ sky130_fd_sc_hd__o31ai_2
X_14007_ _17968_/Q _14036_/A _14006_/Y _14037_/C1 vssd1 vssd1 vccd1 vccd1 _17968_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_269_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11219_ _11219_/A _11219_/B vssd1 vssd1 vccd1 vccd1 _11219_/Y sky130_fd_sc_hd__nor2_1
X_12199_ _17863_/Q _12200_/C _17864_/Q vssd1 vssd1 vccd1 vccd1 _12201_/B sky130_fd_sc_hd__a21oi_1
XFILLER_268_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18815_ _19619_/CLK _18815_/D vssd1 vssd1 vccd1 vccd1 _18815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18746_ _18746_/CLK _18746_/D vssd1 vssd1 vccd1 vccd1 _18746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15958_ _18694_/Q _15970_/A2 _15976_/B1 _18743_/Q _15976_/C1 vssd1 vssd1 vccd1 vccd1
+ _15958_/X sky130_fd_sc_hd__a221o_1
XFILLER_255_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput190 localMemory_wb_adr_i[0] vssd1 vssd1 vccd1 vccd1 input190/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ _14905_/Y _14908_/X _15010_/B1 vssd1 vssd1 vccd1 vccd1 _14909_/Y sky130_fd_sc_hd__a21oi_4
X_18677_ _18683_/CLK _18677_/D vssd1 vssd1 vccd1 vccd1 _18677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15889_ _18672_/Q _15910_/A2 _15888_/X _15904_/C1 vssd1 vssd1 vccd1 vccd1 _18672_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17628_ _17694_/A0 _19556_/Q _17648_/S vssd1 vssd1 vccd1 vccd1 _19556_/D sky130_fd_sc_hd__mux2_1
XFILLER_252_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17559_ _17559_/A _17559_/B vssd1 vssd1 vccd1 vccd1 _17559_/X sky130_fd_sc_hd__and2_1
XFILLER_149_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19229_ _19229_/CLK _19229_/D vssd1 vssd1 vccd1 vccd1 _19229_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09815_ _12601_/B vssd1 vssd1 vccd1 vccd1 _09818_/B sky130_fd_sc_hd__clkinv_2
XFILLER_274_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09746_ _11251_/S _09744_/X _09745_/X vssd1 vssd1 vccd1 vccd1 _09746_/X sky130_fd_sc_hd__o21a_1
XFILLER_274_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09675_/X _09676_/X _10264_/S vssd1 vssd1 vccd1 vccd1 _09677_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11570_ _11084_/S _11569_/X _11570_/B1 vssd1 vssd1 vccd1 vccd1 _11570_/X sky130_fd_sc_hd__o21a_1
XFILLER_168_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10521_ _11602_/C1 _10514_/X _11286_/B1 vssd1 vssd1 vccd1 vccd1 _10521_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13240_ _19306_/Q _12532_/Y _12536_/Y _15920_/A _12505_/Y vssd1 vssd1 vccd1 vccd1
+ _13240_/X sky130_fd_sc_hd__a221o_1
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10452_ _10453_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _13797_/S sky130_fd_sc_hd__and2_2
XFILLER_136_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13171_ _19432_/Q _12560_/B _13169_/X _13170_/X vssd1 vssd1 vccd1 vccd1 _13171_/X
+ sky130_fd_sc_hd__o22a_1
X_10383_ _17978_/Q _11447_/A2 _11371_/B1 vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__a21o_1
XFILLER_272_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12122_ _17835_/Q _12122_/B vssd1 vssd1 vccd1 vccd1 _12128_/C sky130_fd_sc_hd__and2_2
Xclkbuf_leaf_33_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19592_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16930_ _16836_/S _17941_/Q _16929_/X vssd1 vssd1 vccd1 vccd1 _17184_/B sky130_fd_sc_hd__o21a_4
X_12053_ _12053_/A _12073_/B vssd1 vssd1 vccd1 vccd1 _12053_/X sky130_fd_sc_hd__or2_1
XFILLER_111_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1801 _17799_/Q vssd1 vssd1 vccd1 vccd1 _16392_/B sky130_fd_sc_hd__buf_6
XFILLER_284_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1812 _17374_/A vssd1 vssd1 vccd1 vccd1 _15718_/C1 sky130_fd_sc_hd__buf_2
XFILLER_104_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1823 _14342_/A vssd1 vssd1 vccd1 vccd1 _14340_/A sky130_fd_sc_hd__buf_6
XFILLER_78_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11004_ _18457_/Q _18358_/Q _11477_/S vssd1 vssd1 vccd1 vccd1 _11004_/X sky130_fd_sc_hd__mux2_1
Xfanout1834 _14417_/A vssd1 vssd1 vccd1 vccd1 _12383_/C1 sky130_fd_sc_hd__buf_4
X_16861_ _12492_/A _17924_/Q _16860_/X vssd1 vssd1 vccd1 vccd1 _17567_/A sky130_fd_sc_hd__o21a_4
Xfanout1845 _17322_/A vssd1 vssd1 vccd1 vccd1 _17378_/A sky130_fd_sc_hd__buf_4
Xfanout1856 fanout1863/X vssd1 vssd1 vccd1 vccd1 _16153_/D sky130_fd_sc_hd__buf_4
Xfanout1867 _16780_/B1 vssd1 vssd1 vccd1 vccd1 _16764_/B1 sky130_fd_sc_hd__buf_2
XFILLER_237_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout880 _10089_/B vssd1 vssd1 vccd1 vccd1 _15832_/A1 sky130_fd_sc_hd__clkbuf_2
X_18600_ _18632_/CLK _18600_/D vssd1 vssd1 vccd1 vccd1 _18600_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1878 _14423_/B vssd1 vssd1 vccd1 vccd1 _17255_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_266_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1889 _12187_/A vssd1 vssd1 vccd1 vccd1 _12107_/A sky130_fd_sc_hd__buf_4
X_15812_ _18604_/Q _16602_/A0 _15829_/S vssd1 vssd1 vccd1 vccd1 _18604_/D sky130_fd_sc_hd__mux2_1
Xfanout891 _13134_/S vssd1 vssd1 vccd1 vccd1 _13041_/S sky130_fd_sc_hd__buf_2
X_19580_ _19612_/CLK _19580_/D vssd1 vssd1 vccd1 vccd1 _19580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16792_ _16795_/A _16792_/B _16794_/B vssd1 vssd1 vccd1 vccd1 _19285_/D sky130_fd_sc_hd__nor3_1
XFILLER_203_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18531_ _19464_/CLK _18531_/D vssd1 vssd1 vccd1 vccd1 _18531_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_234_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15743_ _18130_/Q _15763_/A2 _15742_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _15744_/B
+ sky130_fd_sc_hd__o22a_2
X_12955_ _13602_/B2 _12947_/X _12954_/X vssd1 vssd1 vccd1 vccd1 _12955_/Y sky130_fd_sc_hd__o21ai_4
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ _14141_/B _11834_/B _11875_/Y vssd1 vssd1 vccd1 vccd1 _11906_/X sky130_fd_sc_hd__a21o_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18462_ _19641_/CLK _18462_/D vssd1 vssd1 vccd1 vccd1 _18462_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_240 _18398_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _19481_/Q _15781_/S _15673_/Y _15717_/B2 vssd1 vssd1 vccd1 vccd1 _15674_/X
+ sky130_fd_sc_hd__o211a_1
X_12886_ _12716_/X _12731_/X _12943_/S vssd1 vssd1 vccd1 vccd1 _13089_/B sky130_fd_sc_hd__mux2_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_251 _19230_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 input220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17413_/A _17423_/B vssd1 vssd1 vccd1 vccd1 _17413_/Y sky130_fd_sc_hd__nand2_1
XFILLER_221_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_273 input238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14625_ _16551_/A0 _18432_/Q _14631_/S vssd1 vssd1 vccd1 vccd1 _18432_/D sky130_fd_sc_hd__mux2_1
X_11837_ _11837_/A _11864_/B vssd1 vssd1 vccd1 vccd1 _11837_/X sky130_fd_sc_hd__or2_4
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_284 _11765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18393_ _19399_/CLK _18393_/D vssd1 vssd1 vccd1 vccd1 _18393_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_295 _08883_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17344_ _17559_/A _17344_/B vssd1 vssd1 vccd1 vccd1 _19469_/D sky130_fd_sc_hd__and2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _14586_/A _14556_/B vssd1 vssd1 vccd1 vccd1 _18386_/D sky130_fd_sc_hd__or2_1
X_11768_ _18586_/Q _11726_/B _11818_/B _11643_/Y vssd1 vssd1 vccd1 vccd1 _11768_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_187_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10719_ _10717_/X _10718_/X _10719_/S vssd1 vssd1 vccd1 vccd1 _10719_/X sky130_fd_sc_hd__mux2_1
X_13507_ _13758_/A _13507_/B vssd1 vssd1 vccd1 vccd1 _13507_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14487_ _14487_/A _14487_/B vssd1 vssd1 vccd1 vccd1 _18339_/D sky130_fd_sc_hd__nor2_1
X_17275_ _18119_/Q _17540_/B1 _17483_/A _17313_/B vssd1 vssd1 vccd1 vccd1 _17275_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_174_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11699_ _18581_/Q _18580_/Q _18579_/Q _18578_/Q vssd1 vssd1 vccd1 vccd1 _11701_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_174_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19014_ _19206_/CLK _19014_/D vssd1 vssd1 vccd1 vccd1 _19014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16226_ _16292_/A0 _18842_/Q _16226_/S vssd1 vssd1 vccd1 vccd1 _18842_/D sky130_fd_sc_hd__mux2_1
X_13438_ _13438_/A _13438_/B vssd1 vssd1 vccd1 vccd1 _13438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16157_ _19424_/Q _17352_/A _15416_/A _16156_/Y _16155_/X vssd1 vssd1 vccd1 vccd1
+ _18777_/D sky130_fd_sc_hd__a41o_1
X_13369_ _15404_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _13369_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15108_ _15108_/A _15108_/B vssd1 vssd1 vccd1 vccd1 _15108_/X sky130_fd_sc_hd__xor2_2
X_16088_ _16096_/A1 _16087_/Y _17725_/C1 vssd1 vssd1 vccd1 vccd1 _18746_/D sky130_fd_sc_hd__a21oi_1
XFILLER_170_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15039_ _15039_/A _15039_/B vssd1 vssd1 vccd1 vccd1 _18528_/D sky130_fd_sc_hd__and2_4
XFILLER_123_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09600_ _19104_/Q _19136_/Q _10717_/S vssd1 vssd1 vccd1 vccd1 _09600_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09531_ _09845_/S _09526_/X _09530_/X vssd1 vssd1 vccd1 vccd1 _09531_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18729_ _18734_/CLK _18729_/D vssd1 vssd1 vccd1 vccd1 _18729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09462_ _18601_/Q _18172_/Q _09464_/S vssd1 vssd1 vccd1 vccd1 _09462_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09393_ _10354_/A1 _18212_/Q _10353_/S _18947_/Q _09381_/S vssd1 vssd1 vccd1 vccd1
+ _09393_/X sky130_fd_sc_hd__o221a_1
XFILLER_178_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput450 _18101_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[0] sky130_fd_sc_hd__buf_4
Xoutput461 _18102_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[1] sky130_fd_sc_hd__buf_4
XFILLER_121_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput472 _18103_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[2] sky130_fd_sc_hd__buf_4
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput483 _11718_/Y vssd1 vssd1 vccd1 vccd1 web0 sky130_fd_sc_hd__buf_4
Xfanout1108 _12587_/Y vssd1 vssd1 vccd1 vccd1 _13930_/A1 sky130_fd_sc_hd__buf_6
Xfanout1119 _12447_/Y vssd1 vssd1 vccd1 vccd1 _13968_/B2 sky130_fd_sc_hd__buf_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire1236 _14417_/B vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__buf_6
XFILLER_219_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09729_ _09978_/A1 _09723_/X _09726_/X _08904_/A vssd1 vssd1 vccd1 vccd1 _09729_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_151_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19530_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12740_ _12740_/A _12740_/B _12740_/C vssd1 vssd1 vccd1 vccd1 _12740_/X sky130_fd_sc_hd__or3_2
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12729_/A _12733_/S vssd1 vssd1 vccd1 vccd1 _12671_/X sky130_fd_sc_hd__or2_1
XFILLER_270_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _17717_/A0 _18261_/Q _14416_/S vssd1 vssd1 vccd1 vccd1 _18261_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11622_ _11622_/A1 _11616_/X _11619_/X _11622_/C1 vssd1 vssd1 vccd1 vccd1 _11622_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15412_/B _15390_/B vssd1 vssd1 vccd1 vccd1 _15390_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14341_ _14341_/A vssd1 vssd1 vccd1 vccd1 _18268_/D sky130_fd_sc_hd__inv_2
XFILLER_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ _11636_/A _11553_/B vssd1 vssd1 vccd1 vccd1 _11635_/A sky130_fd_sc_hd__nand2_2
XFILLER_195_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17060_ _19363_/Q _17113_/B _17059_/Y _16968_/A vssd1 vssd1 vccd1 vccd1 _19363_/D
+ sky130_fd_sc_hd__o211a_1
X_10504_ _10881_/S1 _10493_/X _10503_/X _11621_/C1 vssd1 vssd1 vccd1 vccd1 _10504_/X
+ sky130_fd_sc_hd__o211a_1
X_14272_ _16459_/A _14272_/B vssd1 vssd1 vccd1 vccd1 _17691_/A sky130_fd_sc_hd__nor2_8
X_11484_ _11456_/X _11459_/X _11484_/B1 vssd1 vssd1 vccd1 vccd1 _11484_/X sky130_fd_sc_hd__a21o_1
X_16011_ _18721_/Q _16019_/A2 _16010_/X _16153_/D vssd1 vssd1 vccd1 vccd1 _18721_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13223_ _14340_/A _13223_/B vssd1 vssd1 vccd1 vccd1 _17929_/D sky130_fd_sc_hd__and2_1
X_10435_ _18620_/Q _18191_/Q _11598_/S vssd1 vssd1 vccd1 vccd1 _10435_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13154_ _13316_/B _12836_/Y _13154_/S vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__mux2_2
XFILLER_124_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10366_ _10366_/A1 _18160_/Q _18806_/Q _10370_/S vssd1 vssd1 vccd1 vccd1 _10366_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12105_ _17828_/Q _12106_/C _12104_/Y vssd1 vssd1 vccd1 vccd1 _17828_/D sky130_fd_sc_hd__o21a_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _17982_/CLK _17962_/D vssd1 vssd1 vccd1 vccd1 _17962_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13085_ _13312_/A _14142_/C _13081_/X _13227_/C1 vssd1 vssd1 vccd1 vccd1 _13085_/X
+ sky130_fd_sc_hd__a211o_1
X_10297_ _10297_/A1 _10287_/X _10288_/X vssd1 vssd1 vccd1 vccd1 _10297_/X sky130_fd_sc_hd__o21a_1
XFILLER_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16913_ _18759_/Q _16969_/A2 _16969_/B1 input223/X _16969_/C1 vssd1 vssd1 vccd1 vccd1
+ _16913_/X sky130_fd_sc_hd__a221o_2
Xfanout1620 _09010_/Y vssd1 vssd1 vccd1 vccd1 _09907_/A sky130_fd_sc_hd__clkbuf_4
X_12036_ _17893_/Q _12052_/A2 _12035_/Y _12383_/C1 vssd1 vssd1 vccd1 vccd1 _17795_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1631 _12024_/A vssd1 vssd1 vccd1 vccd1 _09285_/C sky130_fd_sc_hd__buf_12
X_17893_ _17958_/CLK _17893_/D vssd1 vssd1 vccd1 vccd1 _17893_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1642 _10817_/A1 vssd1 vssd1 vccd1 vccd1 _11596_/A1 sky130_fd_sc_hd__buf_6
Xfanout1653 _10282_/A1 vssd1 vssd1 vccd1 vccd1 _11190_/A1 sky130_fd_sc_hd__buf_6
XFILLER_265_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1664 _10144_/B1 vssd1 vssd1 vccd1 vccd1 _10293_/B1 sky130_fd_sc_hd__buf_6
XFILLER_144_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19632_ _19632_/CLK _19632_/D vssd1 vssd1 vccd1 vccd1 _19632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16844_ _09028_/B _15843_/B _16848_/S vssd1 vssd1 vccd1 vccd1 _16846_/B sky130_fd_sc_hd__mux2_2
Xfanout1675 _11312_/A1 vssd1 vssd1 vccd1 vccd1 _11572_/A1 sky130_fd_sc_hd__buf_6
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1686 _10323_/A1 vssd1 vssd1 vccd1 vccd1 _11172_/A1 sky130_fd_sc_hd__buf_6
XFILLER_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1697 _09272_/A1 vssd1 vssd1 vccd1 vccd1 _11458_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_281_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19563_ _19595_/CLK _19563_/D vssd1 vssd1 vccd1 vccd1 _19563_/Q sky130_fd_sc_hd__dfxtp_1
X_16775_ _19279_/Q _19278_/Q _16775_/C vssd1 vssd1 vccd1 vccd1 _16778_/B sky130_fd_sc_hd__and3_1
XFILLER_253_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13987_ _17958_/Q _14004_/A _13986_/Y _13987_/C1 vssd1 vssd1 vccd1 vccd1 _17958_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_280_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18514_ _18517_/CLK _18514_/D vssd1 vssd1 vccd1 vccd1 _18514_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15726_ _15744_/A _15726_/B vssd1 vssd1 vccd1 vccd1 _15726_/Y sky130_fd_sc_hd__nand2_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _12942_/S _12938_/B vssd1 vssd1 vccd1 vccd1 _12938_/Y sky130_fd_sc_hd__nand2_1
X_19494_ _19526_/CLK _19494_/D vssd1 vssd1 vccd1 vccd1 _19494_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18445_ _18445_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15657_ _13770_/Y _15110_/X _10524_/Y _15111_/A vssd1 vssd1 vccd1 vccd1 _15657_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _12869_/A vssd1 vssd1 vccd1 vccd1 _12869_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14608_ _16501_/A0 _18415_/Q _14630_/S vssd1 vssd1 vccd1 vccd1 _18415_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18376_ _19465_/CLK _18376_/D vssd1 vssd1 vccd1 vccd1 _18376_/Q sky130_fd_sc_hd__dfxtp_4
X_15588_ _19477_/Q _19411_/Q vssd1 vssd1 vccd1 vccd1 _15590_/A sky130_fd_sc_hd__and2_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17327_ _19461_/Q _17569_/A _17345_/S vssd1 vssd1 vccd1 vccd1 _17328_/B sky130_fd_sc_hd__mux2_1
XFILLER_175_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14539_ _18378_/Q _14559_/A2 _14559_/B1 input37/X vssd1 vssd1 vccd1 vccd1 _14540_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17258_ _17256_/Y _17257_/X _17159_/A vssd1 vssd1 vccd1 vccd1 _19436_/D sky130_fd_sc_hd__a21oi_1
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16209_ _16606_/A0 _18825_/Q _16226_/S vssd1 vssd1 vccd1 vccd1 _18825_/D sky130_fd_sc_hd__mux2_1
XFILLER_255_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17189_ _17285_/A _17189_/B vssd1 vssd1 vccd1 vccd1 _19414_/D sky130_fd_sc_hd__nor2_1
XFILLER_143_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ _08960_/X _08961_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _08962_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08893_ _11607_/S _12023_/A vssd1 vssd1 vccd1 vccd1 _08893_/Y sky130_fd_sc_hd__nor2_8
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09514_ _18054_/Q _10364_/B _09513_/X _09976_/A1 vssd1 vssd1 vccd1 vccd1 _09514_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _18539_/Q _10249_/S vssd1 vssd1 vccd1 vccd1 _09445_/X sky130_fd_sc_hd__or2_1
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09376_ _09708_/A _09376_/B vssd1 vssd1 vccd1 vccd1 _09376_/Y sky130_fd_sc_hd__nand2_1
XFILLER_197_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10220_ _10217_/X _10218_/X _10219_/X _10297_/A1 _10301_/S vssd1 vssd1 vccd1 vccd1
+ _10220_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ _10149_/X _10150_/X _10225_/S vssd1 vssd1 vccd1 vccd1 _10151_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput291 _11966_/X vssd1 vssd1 vccd1 vccd1 addr0[6] sky130_fd_sc_hd__buf_4
X_10082_ _17982_/Q _11447_/A2 _11371_/B1 vssd1 vssd1 vccd1 vccd1 _10082_/X sky130_fd_sc_hd__a21o_1
XFILLER_248_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13910_ _13938_/B _13958_/B _13909_/Y vssd1 vssd1 vccd1 vccd1 _13910_/X sky130_fd_sc_hd__o21a_1
X_14890_ _18490_/Q _15011_/A2 _14889_/Y _16795_/A vssd1 vssd1 vccd1 vccd1 _18490_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_235_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13841_ _17915_/Q _12448_/C _12762_/B _13840_/Y vssd1 vssd1 vccd1 vccd1 _13841_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_47_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16560_ _16593_/A0 _19164_/Q _16589_/S vssd1 vssd1 vccd1 vccd1 _19164_/D sky130_fd_sc_hd__mux2_1
X_13772_ _13739_/A _13761_/A _13771_/X vssd1 vssd1 vccd1 vccd1 _13772_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10984_ _10984_/A vssd1 vssd1 vccd1 vccd1 _11673_/A sky130_fd_sc_hd__inv_2
XFILLER_204_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15511_ _15511_/A _15511_/B vssd1 vssd1 vccd1 vccd1 _15511_/Y sky130_fd_sc_hd__xnor2_1
X_12723_ _11212_/Y _12595_/B _12729_/B vssd1 vssd1 vccd1 vccd1 _12723_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16491_ _16557_/A0 _19098_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _19098_/D sky130_fd_sc_hd__mux2_1
XFILLER_203_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18230_ _19157_/CLK _18230_/D vssd1 vssd1 vccd1 vccd1 _18230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12654_ _13812_/A _12652_/Y _12653_/Y vssd1 vssd1 vccd1 vccd1 _12654_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15442_ _19471_/Q _19405_/Q vssd1 vssd1 vccd1 vccd1 _15444_/A sky130_fd_sc_hd__nand2_1
XFILLER_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11605_ _19649_/Q _18938_/Q _11605_/S vssd1 vssd1 vccd1 vccd1 _11605_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18161_ _19646_/CLK _18161_/D vssd1 vssd1 vccd1 vccd1 _18161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12585_ _13929_/A1 _12550_/X _12453_/X vssd1 vssd1 vccd1 vccd1 _12585_/X sky130_fd_sc_hd__a21o_1
X_15373_ _15373_/A _15373_/B vssd1 vssd1 vccd1 vccd1 _15376_/A sky130_fd_sc_hd__nand2_2
XFILLER_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17112_ _17208_/B _17116_/A2 _17111_/X _17368_/A vssd1 vssd1 vccd1 vccd1 _19389_/D
+ sky130_fd_sc_hd__o211a_1
X_14324_ _18181_/Q _16542_/A0 _14335_/S vssd1 vssd1 vccd1 vccd1 _18181_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11536_ _11537_/B _13600_/S _10831_/A vssd1 vssd1 vccd1 vccd1 _11536_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18092_ _19306_/CLK _18092_/D vssd1 vssd1 vccd1 vccd1 _18092_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_184_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17043_ _19358_/Q _17043_/B vssd1 vssd1 vccd1 vccd1 _17043_/X sky130_fd_sc_hd__or2_1
X_14255_ _18299_/Q _14261_/A2 _14254_/X _14450_/B vssd1 vssd1 vccd1 vccd1 _18125_/D
+ sky130_fd_sc_hd__o211a_1
X_11467_ _18451_/Q _11477_/S _09129_/S vssd1 vssd1 vccd1 vccd1 _11467_/X sky130_fd_sc_hd__o21a_1
XFILLER_171_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13206_ _19305_/Q _13952_/A2 _12536_/Y _15917_/A _12505_/Y vssd1 vssd1 vccd1 vccd1
+ _13206_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10418_ _18558_/Q _18433_/Q _10426_/S vssd1 vssd1 vccd1 vccd1 _10418_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14186_ _18704_/Q _18091_/Q _14186_/S vssd1 vssd1 vccd1 vccd1 _14187_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11398_ _09099_/A _11393_/X _11397_/X _12466_/A0 vssd1 vssd1 vccd1 vccd1 _11398_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13137_ _13137_/A vssd1 vssd1 vccd1 vccd1 _13137_/Y sky130_fd_sc_hd__inv_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10349_ _18653_/Q _10353_/S vssd1 vssd1 vccd1 vccd1 _10349_/X sky130_fd_sc_hd__or2_1
XFILLER_151_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18994_ _19154_/CLK _18994_/D vssd1 vssd1 vccd1 vccd1 _18994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17945_ _18627_/CLK _17945_/D vssd1 vssd1 vccd1 vccd1 _17945_/Q sky130_fd_sc_hd__dfxtp_2
X_13068_ _19366_/Q _12570_/C _13062_/Y _13067_/X _12570_/D vssd1 vssd1 vccd1 vccd1
+ _13068_/X sky130_fd_sc_hd__a221o_2
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12019_ _17786_/Q _16488_/A0 _12019_/S vssd1 vssd1 vccd1 vccd1 _17786_/D sky130_fd_sc_hd__mux2_1
Xfanout1450 _09857_/A1 vssd1 vssd1 vccd1 vccd1 _11569_/S1 sky130_fd_sc_hd__buf_6
Xfanout1461 _08902_/Y vssd1 vssd1 vccd1 vccd1 _10217_/B sky130_fd_sc_hd__buf_8
XFILLER_238_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17876_ _19324_/CLK _17876_/D vssd1 vssd1 vccd1 vccd1 _17876_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1472 _10511_/S vssd1 vssd1 vccd1 vccd1 _10656_/S sky130_fd_sc_hd__buf_6
XFILLER_94_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1483 fanout1485/X vssd1 vssd1 vccd1 vccd1 _11617_/S sky130_fd_sc_hd__buf_6
X_19615_ _19615_/CLK _19615_/D vssd1 vssd1 vccd1 vccd1 _19615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_266_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1494 fanout1525/X vssd1 vssd1 vccd1 vccd1 _10721_/S sky130_fd_sc_hd__buf_6
X_16827_ _17811_/Q _14675_/B _16836_/S vssd1 vssd1 vccd1 vccd1 _16973_/B sky130_fd_sc_hd__mux2_2
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19546_ _19546_/CLK _19546_/D vssd1 vssd1 vccd1 vccd1 _19546_/Q sky130_fd_sc_hd__dfxtp_1
X_16758_ _19272_/Q _16759_/C _19273_/Q vssd1 vssd1 vccd1 vccd1 _16760_/B sky130_fd_sc_hd__a21oi_1
XFILLER_253_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15709_ _15690_/A _15706_/Y _15708_/Y _15751_/A vssd1 vssd1 vccd1 vccd1 _15709_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_222_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19477_ _19477_/CLK _19477_/D vssd1 vssd1 vccd1 vccd1 _19477_/Q sky130_fd_sc_hd__dfxtp_4
X_16689_ _16740_/A _16695_/C vssd1 vssd1 vccd1 vccd1 _16689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_221_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09230_ _13230_/S _09230_/B vssd1 vssd1 vccd1 vccd1 _13225_/A sky130_fd_sc_hd__nand2b_4
X_18428_ _19575_/CLK _18428_/D vssd1 vssd1 vccd1 vccd1 _18428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09161_ _18143_/Q _18789_/Q _10099_/S vssd1 vssd1 vccd1 vccd1 _09161_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18359_ _19637_/CLK _18359_/D vssd1 vssd1 vccd1 vccd1 _18359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09092_ _09854_/A _12023_/A vssd1 vssd1 vccd1 vccd1 _09092_/Y sky130_fd_sc_hd__nor2_8
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09994_ _09987_/A _09989_/X _09993_/X _11451_/A2 vssd1 vssd1 vccd1 vccd1 _09994_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08945_ _08941_/X _08943_/Y _08940_/X vssd1 vssd1 vccd1 vccd1 _08945_/X sky130_fd_sc_hd__a21o_4
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08876_ _12435_/A _12437_/A _08876_/C vssd1 vssd1 vccd1 vccd1 _12323_/A sky130_fd_sc_hd__or3_4
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09428_ _10366_/A1 _18601_/Q _18172_/Q _09428_/B2 vssd1 vssd1 vccd1 vccd1 _09428_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09359_ _10336_/A _09357_/X _09358_/X _09137_/S vssd1 vssd1 vccd1 vccd1 _09360_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_212_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12370_ _12382_/A _12370_/B vssd1 vssd1 vccd1 vccd1 _12370_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11321_ _11328_/S _11316_/X _11320_/X _11579_/A vssd1 vssd1 vccd1 vccd1 _11321_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ _17798_/Q _14074_/C _16459_/B vssd1 vssd1 vccd1 vccd1 _16359_/A sky130_fd_sc_hd__or3_2
X_11252_ _11248_/X _11251_/X _11252_/S vssd1 vssd1 vccd1 vccd1 _11252_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10203_ _18655_/Q _18077_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _10203_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ _11189_/A _11183_/B vssd1 vssd1 vccd1 vccd1 _11183_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10134_ _10346_/S _10132_/X _10133_/X _10356_/C1 vssd1 vssd1 vccd1 vccd1 _10134_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _18711_/Q _16005_/A2 _15990_/X _14205_/A vssd1 vssd1 vccd1 vccd1 _18711_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17730_ _18630_/Q vssd1 vssd1 vccd1 vccd1 _18630_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_282_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10065_ _12842_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _11653_/A sky130_fd_sc_hd__nor2_2
X_14942_ _17815_/Q _15002_/B vssd1 vssd1 vccd1 vccd1 _14942_/X sky130_fd_sc_hd__or2_1
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17661_ _17661_/A0 _19588_/Q _17681_/S vssd1 vssd1 vccd1 vccd1 _19588_/D sky130_fd_sc_hd__mux2_1
XFILLER_236_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14873_ _14871_/X _14872_/X _14913_/B1 vssd1 vssd1 vccd1 vccd1 _14873_/X sky130_fd_sc_hd__a21o_1
XFILLER_75_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19400_ _19433_/CLK _19400_/D vssd1 vssd1 vccd1 vccd1 _19400_/Q sky130_fd_sc_hd__dfxtp_1
X_16612_ _17712_/A0 _19215_/Q _16618_/S vssd1 vssd1 vccd1 vccd1 _19215_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13824_ _19517_/Q _13947_/A2 _13947_/B1 _13823_/X vssd1 vssd1 vccd1 vccd1 _13824_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17592_ _19488_/Q _17592_/B vssd1 vssd1 vccd1 vccd1 _17592_/X sky130_fd_sc_hd__and2_4
XFILLER_250_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19331_ _19458_/CLK _19331_/D vssd1 vssd1 vccd1 vccd1 _19331_/Q sky130_fd_sc_hd__dfxtp_1
X_16543_ _16543_/A0 _19148_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _19148_/D sky130_fd_sc_hd__mux2_1
XFILLER_245_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13755_ _13747_/B2 _13744_/X _13746_/Y _13754_/Y vssd1 vssd1 vccd1 vccd1 _14024_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_189_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10967_ _18862_/Q _18894_/Q _19054_/Q _19022_/Q _11340_/B2 _11357_/S1 vssd1 vssd1
+ vccd1 vccd1 _10967_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19262_ _19295_/CLK _19262_/D vssd1 vssd1 vccd1 vccd1 _19262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12706_ _13962_/A _13911_/A vssd1 vssd1 vccd1 vccd1 _12743_/A sky130_fd_sc_hd__or2_1
X_16474_ _16507_/A0 _19081_/Q _16491_/S vssd1 vssd1 vccd1 vccd1 _19081_/D sky130_fd_sc_hd__mux2_1
XFILLER_203_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13686_ _19415_/Q _13948_/A2 _13948_/B1 vssd1 vssd1 vccd1 vccd1 _13686_/X sky130_fd_sc_hd__a21o_1
X_10898_ _11606_/S _10897_/X _11623_/A1 vssd1 vssd1 vccd1 vccd1 _10898_/X sky130_fd_sc_hd__a21o_1
X_18213_ _19140_/CLK _18213_/D vssd1 vssd1 vccd1 vccd1 _18213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15425_ _18576_/Q _15447_/B _15424_/X _17469_/C1 vssd1 vssd1 vccd1 vccd1 _18576_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19193_ _19193_/CLK _19193_/D vssd1 vssd1 vccd1 vccd1 _19193_/Q sky130_fd_sc_hd__dfxtp_1
X_12637_ _13597_/A _13597_/B vssd1 vssd1 vccd1 vccd1 _13615_/A sky130_fd_sc_hd__nand2b_1
XFILLER_12_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18144_ _19206_/CLK _18144_/D vssd1 vssd1 vccd1 vccd1 _18144_/Q sky130_fd_sc_hd__dfxtp_1
X_12568_ _12570_/D vssd1 vssd1 vccd1 vccd1 _12568_/Y sky130_fd_sc_hd__inv_2
X_15356_ _17900_/Q _15429_/A2 _15484_/A vssd1 vssd1 vccd1 vccd1 _15361_/A sky130_fd_sc_hd__o21a_1
XFILLER_200_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14307_ _14351_/A _16194_/B vssd1 vssd1 vccd1 vccd1 _14307_/Y sky130_fd_sc_hd__nor2_2
X_11519_ _09141_/A _15357_/A _11490_/X vssd1 vssd1 vccd1 vccd1 _12625_/B sky130_fd_sc_hd__o21ai_4
XFILLER_117_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18075_ _19596_/CLK _18075_/D vssd1 vssd1 vccd1 vccd1 _18075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12499_ _12499_/A _12513_/B _12538_/A _12528_/C vssd1 vssd1 vccd1 vccd1 _12582_/A
+ sky130_fd_sc_hd__or4_4
X_15287_ _17917_/Q _15369_/A vssd1 vssd1 vccd1 vccd1 _15289_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17026_ _17184_/B _17032_/A2 _17025_/X _17360_/A vssd1 vssd1 vccd1 vccd1 _19349_/D
+ sky130_fd_sc_hd__o211a_1
X_14238_ _14238_/A _14266_/B vssd1 vssd1 vccd1 vccd1 _14238_/X sky130_fd_sc_hd__or2_1
XFILLER_259_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ _16892_/A _14169_/B vssd1 vssd1 vccd1 vccd1 _18082_/D sky130_fd_sc_hd__and2_1
XFILLER_140_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout709 _13115_/C1 vssd1 vssd1 vccd1 vccd1 _13722_/B1 sky130_fd_sc_hd__buf_8
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18977_ _19147_/CLK _18977_/D vssd1 vssd1 vccd1 vccd1 _18977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _17930_/CLK _17928_/D vssd1 vssd1 vccd1 vccd1 _17928_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_285_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1280 _15970_/A2 vssd1 vssd1 vccd1 vccd1 _15953_/B sky130_fd_sc_hd__buf_4
XFILLER_66_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1291 _14591_/B1 vssd1 vssd1 vccd1 vccd1 _14559_/B1 sky130_fd_sc_hd__buf_4
X_17859_ _18691_/CLK _17859_/D vssd1 vssd1 vccd1 vccd1 _17859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19529_ _19533_/CLK _19529_/D vssd1 vssd1 vccd1 vccd1 _19529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ _10219_/A1 _19564_/Q _10353_/S _19596_/Q _10205_/S vssd1 vssd1 vccd1 vccd1
+ _09213_/X sky130_fd_sc_hd__o221a_1
XFILLER_22_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09144_ _11490_/B _15332_/A _09144_/C vssd1 vssd1 vccd1 vccd1 _13267_/A sky130_fd_sc_hd__and3_2
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09075_ _15307_/A _15082_/A _12443_/B vssd1 vssd1 vccd1 vccd1 _09075_/X sky130_fd_sc_hd__or3_2
XFILLER_135_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09977_ _09978_/A1 _09967_/X _09976_/X _11516_/B1 vssd1 vssd1 vccd1 vccd1 _09977_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ _17796_/Q _17794_/Q vssd1 vssd1 vccd1 vccd1 _08929_/D sky130_fd_sc_hd__nand2_1
XFILLER_58_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08859_ _16787_/A vssd1 vssd1 vccd1 vccd1 _08859_/Y sky130_fd_sc_hd__inv_2
XFILLER_218_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_58_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19613_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _14141_/B _11834_/B _11859_/B vssd1 vssd1 vccd1 vccd1 _11870_/X sky130_fd_sc_hd__o21a_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _19639_/Q _18928_/Q _11598_/S vssd1 vssd1 vccd1 vccd1 _10821_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ _10753_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _10754_/A sky130_fd_sc_hd__and2_4
XFILLER_38_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13540_ _18119_/Q _13541_/B vssd1 vssd1 vccd1 vccd1 _13606_/C sky130_fd_sc_hd__and2_2
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13471_ _13464_/Y _13467_/Y _13470_/X _13966_/C1 vssd1 vssd1 vccd1 vccd1 _13471_/X
+ sky130_fd_sc_hd__a22o_1
X_10683_ _18461_/Q _18362_/Q _11249_/S vssd1 vssd1 vccd1 vccd1 _10683_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12422_ _17915_/Q _12421_/A _12421_/Y _12428_/C1 vssd1 vssd1 vccd1 vccd1 _17915_/D
+ sky130_fd_sc_hd__o211a_1
X_15210_ _19429_/Q _15411_/B _17151_/A _15209_/X vssd1 vssd1 vccd1 vccd1 _15210_/X
+ sky130_fd_sc_hd__o211a_1
X_16190_ _16455_/A1 _18807_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _18807_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12353_ _17892_/Q _12349_/A _12352_/Y _12383_/C1 vssd1 vssd1 vccd1 vccd1 _17892_/D
+ sky130_fd_sc_hd__o211a_1
X_15141_ _19457_/Q _17559_/B _19456_/Q vssd1 vssd1 vccd1 vccd1 _15523_/S sky130_fd_sc_hd__nor3b_4
XFILLER_127_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11304_ _11305_/A1 _18218_/Q _11309_/S _18953_/Q _11311_/C1 vssd1 vssd1 vccd1 vccd1
+ _11304_/X sky130_fd_sc_hd__o221a_1
X_15072_ _18556_/Q _17683_/A0 _15079_/S vssd1 vssd1 vccd1 vccd1 _18556_/D sky130_fd_sc_hd__mux2_1
X_12284_ _12474_/B _12483_/B _12476_/B vssd1 vssd1 vccd1 vccd1 _12284_/X sky130_fd_sc_hd__and3_1
X_14023_ _14033_/A1 _13723_/X _14022_/X _14179_/A vssd1 vssd1 vccd1 vccd1 _17976_/D
+ sky130_fd_sc_hd__o211a_1
X_18900_ _19643_/CLK _18900_/D vssd1 vssd1 vccd1 vccd1 _18900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11235_ _11250_/A1 _19569_/Q _11247_/S _19601_/Q _11569_/S1 vssd1 vssd1 vccd1 vccd1
+ _11235_/X sky130_fd_sc_hd__o221a_1
XFILLER_268_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18831_ _19575_/CLK _18831_/D vssd1 vssd1 vccd1 vccd1 _18831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11166_ _10689_/S _11161_/X _11165_/X _08843_/A vssd1 vssd1 vccd1 vccd1 _11166_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10117_ _10250_/S _10116_/X _11459_/B1 vssd1 vssd1 vccd1 vccd1 _10117_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18762_ _18772_/CLK _18762_/D vssd1 vssd1 vccd1 vccd1 _18762_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_209_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15974_ _18702_/Q _15953_/B _16002_/B1 _18751_/Q _16002_/C1 vssd1 vssd1 vccd1 vccd1
+ _15974_/X sky130_fd_sc_hd__a221o_1
X_11097_ _11091_/X _11093_/X _11096_/X _11578_/S _11588_/B1 vssd1 vssd1 vccd1 vccd1
+ _11097_/X sky130_fd_sc_hd__o221a_1
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _17713_/A0 _19639_/Q _17718_/S vssd1 vssd1 vccd1 vccd1 _19639_/D sky130_fd_sc_hd__mux2_1
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14925_ _15006_/A1 _14924_/X _15006_/B1 vssd1 vssd1 vccd1 vccd1 _14925_/Y sky130_fd_sc_hd__o21ai_2
X_10048_ _11618_/A1 _19554_/Q _10726_/S _19586_/Q _10745_/S vssd1 vssd1 vccd1 vccd1
+ _10048_/X sky130_fd_sc_hd__o221a_1
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18693_ _18738_/CLK _18693_/D vssd1 vssd1 vccd1 vccd1 _18693_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17644_ _17644_/A0 _19572_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _19572_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856_ input50/X input85/X _14947_/S vssd1 vssd1 vccd1 vccd1 _14857_/A sky130_fd_sc_hd__mux2_2
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13807_ _13807_/A _13807_/B vssd1 vssd1 vccd1 vccd1 _13807_/X sky130_fd_sc_hd__or2_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17575_ _17575_/A _17589_/B vssd1 vssd1 vccd1 vccd1 _17575_/X sky130_fd_sc_hd__or2_1
X_14787_ _14783_/Y _14786_/X _14879_/B1 vssd1 vssd1 vccd1 vccd1 _14787_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11999_ _17766_/Q _16501_/A0 _12021_/S vssd1 vssd1 vccd1 vccd1 _17766_/D sky130_fd_sc_hd__mux2_1
X_19314_ _19326_/CLK _19314_/D vssd1 vssd1 vccd1 vccd1 _19314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16526_ _16526_/A0 _19131_/Q _16548_/S vssd1 vssd1 vccd1 vccd1 _19131_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13738_ _15133_/A _13734_/X _13737_/X _13869_/B2 vssd1 vssd1 vccd1 vccd1 _13739_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19245_ _19280_/CLK _19245_/D vssd1 vssd1 vccd1 vccd1 _19245_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_231_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16457_ _19065_/Q _16490_/A0 _16457_/S vssd1 vssd1 vccd1 vccd1 _19065_/D sky130_fd_sc_hd__mux2_1
X_13669_ _13896_/B2 _13197_/X _13668_/X _13966_/C1 vssd1 vssd1 vccd1 vccd1 _13669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15408_ _15408_/A _15408_/B vssd1 vssd1 vccd1 vccd1 _15456_/C sky130_fd_sc_hd__xnor2_4
X_19176_ _19208_/CLK _19176_/D vssd1 vssd1 vccd1 vccd1 _19176_/Q sky130_fd_sc_hd__dfxtp_1
X_16388_ _16488_/A0 _18999_/Q _16388_/S vssd1 vssd1 vccd1 vccd1 _18999_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18127_ _19453_/CLK _18127_/D vssd1 vssd1 vccd1 vccd1 _18127_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15339_ _15308_/B _15313_/B _15365_/D _15307_/B vssd1 vssd1 vccd1 vccd1 _15340_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_247_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18058_ _19636_/CLK _18058_/D vssd1 vssd1 vccd1 vccd1 _18058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09900_ _17953_/Q _11447_/A2 _11371_/B1 vssd1 vssd1 vccd1 vccd1 _09900_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_172_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17009_ _19341_/Q _17009_/B vssd1 vssd1 vccd1 vccd1 _17009_/X sky130_fd_sc_hd__or2_1
XFILLER_104_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout506 _17523_/B vssd1 vssd1 vccd1 vccd1 _17493_/B sky130_fd_sc_hd__buf_4
XFILLER_263_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout517 _17244_/B vssd1 vssd1 vccd1 vccd1 _17310_/B sky130_fd_sc_hd__buf_4
X_09831_ _18238_/Q _10001_/S _10707_/A _09830_/X vssd1 vssd1 vccd1 vccd1 _09831_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout528 _11770_/B1 vssd1 vssd1 vccd1 vccd1 _11844_/A sky130_fd_sc_hd__buf_4
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout539 _15633_/C1 vssd1 vssd1 vccd1 vccd1 _15499_/B1 sky130_fd_sc_hd__buf_4
XFILLER_101_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09762_ _11565_/A1 _19134_/Q _11070_/S _19102_/Q vssd1 vssd1 vccd1 vccd1 _09762_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_258_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09693_ _09611_/A _09692_/X _11790_/B vssd1 vssd1 vccd1 vccd1 _09693_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_39_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_176_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19444_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09127_ _09125_/X _09126_/X _09264_/S vssd1 vssd1 vccd1 vccd1 _09127_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_105_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18713_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_135_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09058_ _12598_/A vssd1 vssd1 vccd1 vccd1 _09143_/A sky130_fd_sc_hd__clkinv_2
XFILLER_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11020_ _10993_/X _10996_/X _11484_/B1 vssd1 vssd1 vccd1 vccd1 _11020_/X sky130_fd_sc_hd__a21o_1
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _19428_/Q _12560_/B _12969_/X _12970_/X _12560_/A vssd1 vssd1 vccd1 vccd1
+ _12971_/X sky130_fd_sc_hd__o221a_1
XFILLER_218_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _14720_/A _14710_/B vssd1 vssd1 vccd1 vccd1 _14710_/Y sky130_fd_sc_hd__nor2_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11926_/A1 _11939_/A1 _11846_/B _11935_/B1 input237/X vssd1 vssd1 vccd1 vccd1
+ _11922_/X sky130_fd_sc_hd__a32o_4
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15690_ _15690_/A _15690_/B vssd1 vssd1 vccd1 vccd1 _15690_/Y sky130_fd_sc_hd__nor2_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_400 _12609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_411 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_422 _12956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14641_ _17700_/A0 _18447_/Q _14660_/S vssd1 vssd1 vccd1 vccd1 _18447_/D sky130_fd_sc_hd__mux2_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_433 _11904_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_444 _13477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11853_ _11909_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11853_/X sky130_fd_sc_hd__and2_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_455 _18573_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_466 _18374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_477 input227/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ _19088_/Q _18992_/Q _11605_/S vssd1 vssd1 vccd1 vccd1 _10804_/X sky130_fd_sc_hd__mux2_1
X_17360_ _17360_/A _17360_/B vssd1 vssd1 vccd1 vccd1 _19477_/D sky130_fd_sc_hd__and2_1
XFILLER_25_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_488 _18111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11784_ _11799_/A _11799_/B _11803_/B vssd1 vssd1 vccd1 vccd1 _11784_/X sky130_fd_sc_hd__and3_1
XFILLER_82_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14572_ _14576_/A _14572_/B vssd1 vssd1 vccd1 vccd1 _18394_/D sky130_fd_sc_hd__or2_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_499 _14660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16311_ _17709_/A0 _18924_/Q _16325_/S vssd1 vssd1 vccd1 vccd1 _18924_/D sky130_fd_sc_hd__mux2_1
X_13523_ _19442_/Q _13655_/A2 _13521_/X _13522_/X _13655_/C1 vssd1 vssd1 vccd1 vccd1
+ _13523_/X sky130_fd_sc_hd__o221a_1
X_10735_ _11277_/A1 _19217_/Q _19185_/Q _10370_/S _12766_/A0 vssd1 vssd1 vccd1 vccd1
+ _10735_/X sky130_fd_sc_hd__a221o_1
X_17291_ _17289_/Y _17290_/X _17198_/A vssd1 vssd1 vccd1 vccd1 _19447_/D sky130_fd_sc_hd__a21oi_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19030_ _19623_/CLK _19030_/D vssd1 vssd1 vccd1 vccd1 _19030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16242_ _16606_/A0 _18857_/Q _16259_/S vssd1 vssd1 vccd1 vccd1 _18857_/D sky130_fd_sc_hd__mux2_1
X_10666_ _18462_/Q _18363_/Q _10667_/S vssd1 vssd1 vccd1 vccd1 _10666_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13454_ _19440_/Q _13655_/A2 _13452_/X _13453_/X _13655_/C1 vssd1 vssd1 vccd1 vccd1
+ _13454_/X sky130_fd_sc_hd__o221a_1
XFILLER_185_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12405_ _12429_/A1 _09236_/A _09486_/X _12429_/B1 _18395_/Q vssd1 vssd1 vccd1 vccd1
+ _12406_/B sky130_fd_sc_hd__o32ai_2
XFILLER_127_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16173_ _09105_/A _18790_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _18790_/D sky130_fd_sc_hd__mux2_1
X_13385_ _13402_/B _13961_/A vssd1 vssd1 vccd1 vccd1 _13385_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10597_ _11279_/B1 _10580_/X _10595_/X _10596_/Y vssd1 vssd1 vccd1 vccd1 _10597_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15124_ _15330_/A _15124_/B _15124_/C vssd1 vssd1 vccd1 vccd1 _15124_/X sky130_fd_sc_hd__and3_4
X_12336_ _12312_/X _12761_/B _15416_/A _12335_/X _17724_/B vssd1 vssd1 vccd1 vccd1
+ _12336_/X sky130_fd_sc_hd__o41a_1
XFILLER_217_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15055_ _18539_/Q _16500_/A0 _15076_/S vssd1 vssd1 vccd1 vccd1 _18539_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12267_ _12267_/A _12267_/B vssd1 vssd1 vccd1 vccd1 _12314_/B sky130_fd_sc_hd__or2_4
XFILLER_107_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14006_ _14036_/A _14006_/B vssd1 vssd1 vccd1 vccd1 _14006_/Y sky130_fd_sc_hd__nand2_1
X_11218_ _11218_/A _11218_/B vssd1 vssd1 vccd1 vccd1 _11219_/B sky130_fd_sc_hd__nor2_1
X_12198_ _17863_/Q _12200_/C _12197_/Y vssd1 vssd1 vccd1 vccd1 _17863_/D sky130_fd_sc_hd__o21a_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11149_ _11172_/A1 _18220_/Q _11160_/S _18955_/Q _11156_/C1 vssd1 vssd1 vccd1 vccd1
+ _11149_/X sky130_fd_sc_hd__o221a_1
XFILLER_1_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18814_ _19621_/CLK _18814_/D vssd1 vssd1 vccd1 vccd1 _18814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18745_ _19304_/CLK _18745_/D vssd1 vssd1 vccd1 vccd1 _18745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15957_ _18694_/Q _15977_/A2 _15956_/X _14181_/A vssd1 vssd1 vccd1 vccd1 _18694_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput180 irq[3] vssd1 vssd1 vccd1 vccd1 _15092_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_236_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput191 localMemory_wb_adr_i[10] vssd1 vssd1 vccd1 vccd1 input191/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14908_ _14979_/A1 _18271_/Q _14907_/Y _14918_/B1 vssd1 vssd1 vccd1 vccd1 _14908_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_64_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18676_ _18683_/CLK _18676_/D vssd1 vssd1 vccd1 vccd1 _18676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15888_ _18671_/Q _15906_/A2 _15945_/C1 _15887_/X vssd1 vssd1 vccd1 vccd1 _15888_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17627_ _17660_/A0 _19555_/Q _17654_/S vssd1 vssd1 vccd1 vccd1 _19555_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14839_ _17805_/Q _15002_/B vssd1 vssd1 vccd1 vccd1 _14839_/X sky130_fd_sc_hd__or2_1
XFILLER_251_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17558_ _19522_/Q _17558_/B vssd1 vssd1 vccd1 vccd1 _17558_/X sky130_fd_sc_hd__or2_1
XFILLER_205_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_3_wb_clk_i _19652_/A vssd1 vssd1 vccd1 vccd1 _19573_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16509_ _16542_/A0 _19115_/Q _16515_/S vssd1 vssd1 vccd1 vccd1 _19115_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17489_ _19509_/Q _17493_/B _17487_/X _17488_/Y _17356_/A vssd1 vssd1 vccd1 vccd1
+ _19509_/D sky130_fd_sc_hd__o221a_1
X_19228_ _19229_/CLK _19228_/D vssd1 vssd1 vccd1 vccd1 _19228_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_192_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19159_ _19159_/CLK _19159_/D vssd1 vssd1 vccd1 vccd1 _19159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09814_ _09948_/B _15151_/A _09780_/X vssd1 vssd1 vccd1 vccd1 _12601_/B sky130_fd_sc_hd__a21boi_4
XFILLER_87_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09745_ _11565_/A1 _18136_/Q _18782_/Q _09770_/S _09095_/A vssd1 vssd1 vccd1 vccd1
+ _09745_/X sky130_fd_sc_hd__a221o_1
XFILLER_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _11172_/A1 _17762_/Q _09680_/B1 _18311_/Q vssd1 vssd1 vccd1 vccd1 _09676_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_255_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10520_ _12320_/B _10519_/Y _10518_/Y _11602_/C1 vssd1 vssd1 vccd1 vccd1 _10520_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_52_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10451_ _18127_/Q _10450_/Y _13739_/A vssd1 vssd1 vccd1 vccd1 _12648_/B sky130_fd_sc_hd__mux2_4
XFILLER_182_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13170_ _19400_/Q _12570_/A _13244_/B1 vssd1 vssd1 vccd1 vccd1 _13170_/X sky130_fd_sc_hd__a21o_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10382_ _09574_/A _10085_/B _09148_/X _11143_/A1 vssd1 vssd1 vccd1 vccd1 _10382_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ _16811_/A _12121_/B _12122_/B vssd1 vssd1 vccd1 vccd1 _17834_/D sky130_fd_sc_hd__nor3_1
XFILLER_163_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12052_ _17901_/Q _12052_/A2 _12051_/X _13257_/A vssd1 vssd1 vccd1 vccd1 _17803_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1802 _14427_/B vssd1 vssd1 vccd1 vccd1 _16046_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11003_ _09129_/S _11001_/X _11002_/X _11466_/B1 vssd1 vssd1 vccd1 vccd1 _11003_/X
+ sky130_fd_sc_hd__o31a_1
Xfanout1813 _17380_/A vssd1 vssd1 vccd1 vccd1 _17374_/A sky130_fd_sc_hd__buf_2
Xfanout1824 fanout1870/X vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__buf_6
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19629_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16860_ _18746_/Q _12276_/A _16877_/B1 input241/X _12488_/A vssd1 vssd1 vccd1 vccd1
+ _16860_/X sky130_fd_sc_hd__a221o_1
Xfanout1835 _14417_/A vssd1 vssd1 vccd1 vccd1 _12350_/C1 sky130_fd_sc_hd__buf_2
XFILLER_277_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1846 _13987_/C1 vssd1 vssd1 vccd1 vccd1 _17322_/A sky130_fd_sc_hd__buf_4
Xfanout1857 fanout1863/X vssd1 vssd1 vccd1 vccd1 _14197_/A sky130_fd_sc_hd__buf_4
Xfanout870 _10239_/B vssd1 vssd1 vccd1 vccd1 _16455_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1868 _16812_/B1 vssd1 vssd1 vccd1 vccd1 _16780_/B1 sky130_fd_sc_hd__clkbuf_4
X_15811_ _18603_/Q _17701_/A0 _15832_/S vssd1 vssd1 vccd1 vccd1 _18603_/D sky130_fd_sc_hd__mux2_1
XFILLER_265_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout881 _12823_/A vssd1 vssd1 vccd1 vccd1 _12821_/A sky130_fd_sc_hd__buf_4
Xfanout1879 _14487_/A vssd1 vssd1 vccd1 vccd1 _14423_/B sky130_fd_sc_hd__buf_12
X_16791_ _19285_/Q _19284_/Q _16791_/C vssd1 vssd1 vccd1 vccd1 _16794_/B sky130_fd_sc_hd__and3_1
Xfanout892 _09898_/A vssd1 vssd1 vccd1 vccd1 _13134_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_253_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18530_ _19229_/CLK _18530_/D vssd1 vssd1 vccd1 vccd1 _18530_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_234_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15742_ _13874_/A _15502_/B _13903_/B _15112_/B vssd1 vssd1 vccd1 vccd1 _15742_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12954_ _12704_/S _12953_/X _12949_/X _12265_/Y vssd1 vssd1 vccd1 vccd1 _12954_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_206_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _19025_/CLK _18461_/D vssd1 vssd1 vccd1 vccd1 _18461_/Q sky130_fd_sc_hd__dfxtp_1
X_11905_ _11591_/X _11869_/B _11801_/A vssd1 vssd1 vccd1 vccd1 _11908_/A sky130_fd_sc_hd__a21oi_4
XFILLER_206_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _15716_/S _15673_/B vssd1 vssd1 vccd1 vccd1 _15673_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _18390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12885_ _12885_/A vssd1 vssd1 vccd1 vccd1 _12885_/Y sky130_fd_sc_hd__inv_2
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_241 _18398_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_252 _19230_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _18105_/Q _17437_/A2 _17410_/X _17411_/X vssd1 vssd1 vccd1 vccd1 _17412_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_263 input221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14624_ _17683_/A0 _18431_/Q _14631_/S vssd1 vssd1 vccd1 vccd1 _18431_/D sky130_fd_sc_hd__mux2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _11844_/A _11836_/B vssd1 vssd1 vccd1 vccd1 _11836_/X sky130_fd_sc_hd__and2_1
X_18392_ _19465_/CLK _18392_/D vssd1 vssd1 vccd1 vccd1 _18392_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 input239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 _11886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_296 _18733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _19469_/Q _17585_/A _17377_/S vssd1 vssd1 vccd1 vccd1 _17344_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ _18386_/Q _14559_/A2 _14559_/B1 input14/X vssd1 vssd1 vccd1 vccd1 _14556_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_198_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _18585_/Q _14349_/B _11769_/B1 _11668_/Y vssd1 vssd1 vccd1 vccd1 _11767_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13506_ _13637_/A _14008_/B vssd1 vssd1 vccd1 vccd1 _13506_/X sky130_fd_sc_hd__or2_1
X_10718_ _18554_/Q _18429_/Q _10744_/S vssd1 vssd1 vccd1 vccd1 _10718_/X sky130_fd_sc_hd__mux2_1
X_17274_ _19442_/Q _17313_/B vssd1 vssd1 vccd1 vccd1 _17274_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14486_ _18338_/Q _17690_/A0 _14486_/S vssd1 vssd1 vccd1 vccd1 _18338_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11698_ _18577_/Q _18576_/Q _18575_/Q _18574_/Q vssd1 vssd1 vccd1 vccd1 _11701_/B
+ sky130_fd_sc_hd__or4_2
X_19013_ _19203_/CLK _19013_/D vssd1 vssd1 vccd1 vccd1 _19013_/Q sky130_fd_sc_hd__dfxtp_1
X_16225_ _16622_/A0 _18841_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _18841_/D sky130_fd_sc_hd__mux2_1
X_13437_ _13757_/A _14004_/B vssd1 vssd1 vccd1 vccd1 _13437_/X sky130_fd_sc_hd__or2_1
X_10649_ _10649_/A1 _10648_/X _10647_/X _10881_/S1 vssd1 vssd1 vccd1 vccd1 _10649_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16156_ _17219_/A _16156_/B vssd1 vssd1 vccd1 vccd1 _16156_/Y sky130_fd_sc_hd__nor2_1
X_13368_ _17933_/Q _13742_/A2 _13367_/X _14181_/A vssd1 vssd1 vccd1 vccd1 _17933_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15107_ _09980_/Y _12790_/A _15259_/B vssd1 vssd1 vccd1 vccd1 _15108_/B sky130_fd_sc_hd__mux2_4
XFILLER_170_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12319_ _15133_/A _15111_/A vssd1 vssd1 vccd1 vccd1 _12319_/Y sky130_fd_sc_hd__nand2_1
X_16087_ _18746_/Q _16093_/B vssd1 vssd1 vccd1 vccd1 _16087_/Y sky130_fd_sc_hd__nand2_1
X_13299_ _19404_/Q _12579_/Y _12771_/X _13298_/X _12581_/Y vssd1 vssd1 vccd1 vccd1
+ _13299_/X sky130_fd_sc_hd__a221o_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15038_ _18527_/Q input205/X _15038_/S vssd1 vssd1 vccd1 vccd1 _18527_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16989_ _17565_/B _17043_/B vssd1 vssd1 vccd1 vccd1 _16989_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09530_ _09683_/A _09529_/X _10260_/B1 vssd1 vssd1 vccd1 vccd1 _09530_/X sky130_fd_sc_hd__o21a_1
XFILLER_237_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18728_ _18734_/CLK _18728_/D vssd1 vssd1 vccd1 vccd1 _18728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09461_ _18243_/Q _18818_/Q _09464_/S vssd1 vssd1 vccd1 vccd1 _09461_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18659_ _18660_/CLK _18659_/D vssd1 vssd1 vccd1 vccd1 _18659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09392_ _19075_/Q _18979_/Q _10128_/B vssd1 vssd1 vccd1 vccd1 _09392_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput440 _18479_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[8] sky130_fd_sc_hd__buf_4
XFILLER_161_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput451 _18111_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[10] sky130_fd_sc_hd__buf_4
XFILLER_154_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput462 _18121_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[20] sky130_fd_sc_hd__buf_4
Xoutput473 _18131_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[30] sky130_fd_sc_hd__buf_4
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput484 _11953_/X vssd1 vssd1 vccd1 vccd1 wmask0[0] sky130_fd_sc_hd__buf_4
XFILLER_120_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1109 _13758_/A vssd1 vssd1 vccd1 vccd1 _13438_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_248_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09728_ _11199_/S1 _09718_/X _09727_/X _11516_/B1 vssd1 vssd1 vccd1 vccd1 _09728_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_262_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09659_ _09027_/A _09034_/B _09658_/X _10234_/B _09483_/Y vssd1 vssd1 vccd1 vccd1
+ _09660_/C sky130_fd_sc_hd__a32o_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12669_/X _12668_/X _12821_/A vssd1 vssd1 vccd1 vccd1 _12670_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_191_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19643_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11622_/A1 _11611_/X _11620_/X _11621_/C1 vssd1 vssd1 vccd1 vccd1 _11621_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_120_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19300_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14340_ _14340_/A _14345_/B vssd1 vssd1 vccd1 vccd1 _14341_/A sky130_fd_sc_hd__nand2_1
X_11552_ _13794_/A _11639_/B _13812_/A _11549_/X _10308_/A vssd1 vssd1 vccd1 vccd1
+ _11553_/B sky130_fd_sc_hd__a311o_2
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10503_ _10643_/S _10495_/X _10494_/X _10653_/C1 vssd1 vssd1 vccd1 vccd1 _10503_/X
+ sky130_fd_sc_hd__a211o_1
X_11483_ _09099_/A _11478_/X _11480_/X _11482_/X _08843_/Y vssd1 vssd1 vccd1 vccd1
+ _11483_/Y sky130_fd_sc_hd__o221ai_4
X_14271_ _17797_/Q _14272_/B vssd1 vssd1 vccd1 vccd1 _16326_/A sky130_fd_sc_hd__or2_4
XFILLER_155_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ _18720_/Q _15953_/B _16147_/A2 _18769_/Q _16018_/C1 vssd1 vssd1 vccd1 vccd1
+ _16010_/X sky130_fd_sc_hd__a221o_1
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10434_ _18262_/Q _18837_/Q _11598_/S vssd1 vssd1 vccd1 vccd1 _10434_/X sky130_fd_sc_hd__mux2_1
X_13222_ _09281_/Y _13292_/A2 _13221_/Y _13256_/B1 _17929_/Q vssd1 vssd1 vccd1 vccd1
+ _13223_/B sky130_fd_sc_hd__a32o_1
XFILLER_171_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10365_ _18870_/Q _10370_/S _12766_/A0 vssd1 vssd1 vccd1 vccd1 _10365_/X sky130_fd_sc_hd__o21a_1
X_13153_ _13139_/Y _13152_/Y _13194_/S vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__mux2_2
XFILLER_152_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12104_ _12107_/A _12104_/B vssd1 vssd1 vccd1 vccd1 _12104_/Y sky130_fd_sc_hd__nor2_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17961_ _18627_/CLK _17961_/D vssd1 vssd1 vccd1 vccd1 _17961_/Q sky130_fd_sc_hd__dfxtp_1
X_13084_ _13126_/B _13084_/B vssd1 vssd1 vccd1 vccd1 _14142_/C sky130_fd_sc_hd__and2_1
X_10296_ _09708_/A _10291_/X _10295_/X _08895_/A vssd1 vssd1 vccd1 vccd1 _10296_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1610 _16095_/B vssd1 vssd1 vccd1 vccd1 _16093_/B sky130_fd_sc_hd__buf_6
X_16912_ _16960_/A _16912_/B vssd1 vssd1 vccd1 vccd1 _19312_/D sky130_fd_sc_hd__and2_1
X_12035_ _14741_/A _12035_/B vssd1 vssd1 vccd1 vccd1 _12035_/Y sky130_fd_sc_hd__nand2_1
Xfanout1621 _12409_/A2 vssd1 vssd1 vccd1 vccd1 _09236_/A sky130_fd_sc_hd__buf_6
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17892_ _17901_/CLK _17892_/D vssd1 vssd1 vccd1 vccd1 _17892_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_214_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1632 _08865_/Y vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_266_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1643 _11594_/A1 vssd1 vssd1 vccd1 vccd1 _11352_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_77_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1654 _10282_/A1 vssd1 vssd1 vccd1 vccd1 _11497_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_77_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19631_ _19631_/CLK _19631_/D vssd1 vssd1 vccd1 vccd1 _19631_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1665 _10030_/C1 vssd1 vssd1 vccd1 vccd1 _10144_/B1 sky130_fd_sc_hd__buf_6
X_16843_ _17052_/A _17052_/B _16843_/C _16843_/D vssd1 vssd1 vccd1 vccd1 _16843_/X
+ sky130_fd_sc_hd__and4b_4
Xfanout1676 _11584_/A1 vssd1 vssd1 vccd1 vccd1 _11312_/A1 sky130_fd_sc_hd__buf_6
XFILLER_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1687 _12468_/B vssd1 vssd1 vccd1 vccd1 _10323_/A1 sky130_fd_sc_hd__buf_6
XFILLER_265_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1698 _08845_/Y vssd1 vssd1 vccd1 vccd1 _09272_/A1 sky130_fd_sc_hd__buf_4
XFILLER_219_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19562_ _19594_/CLK _19562_/D vssd1 vssd1 vccd1 vccd1 _19562_/Q sky130_fd_sc_hd__dfxtp_1
X_16774_ _19278_/Q _16775_/C _19279_/Q vssd1 vssd1 vccd1 vccd1 _16776_/B sky130_fd_sc_hd__a21oi_1
X_13986_ _14004_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_253_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18513_ _19321_/CLK _18513_/D vssd1 vssd1 vccd1 vccd1 _18513_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15725_ _15725_/A _15725_/B _15702_/B vssd1 vssd1 vccd1 vccd1 _15726_/B sky130_fd_sc_hd__or3b_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12937_ _13046_/A1 _13263_/B _12932_/X vssd1 vssd1 vccd1 vccd1 _12937_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_46_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19493_ _19552_/CLK _19493_/D vssd1 vssd1 vccd1 vccd1 _19493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ _19653_/A _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15656_ _18586_/Q _15718_/A2 _15648_/Y _15655_/X _15718_/C1 vssd1 vssd1 vccd1 vccd1
+ _18586_/D sky130_fd_sc_hd__o221a_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _18103_/Q _12868_/B vssd1 vssd1 vccd1 vccd1 _12869_/A sky130_fd_sc_hd__xnor2_2
XFILLER_261_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14607_ _16500_/A0 _18414_/Q _14628_/S vssd1 vssd1 vccd1 vccd1 _18414_/D sky130_fd_sc_hd__mux2_1
X_18375_ _19483_/CLK _18375_/D vssd1 vssd1 vccd1 vccd1 _18375_/Q sky130_fd_sc_hd__dfxtp_4
X_11819_ _11819_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11819_/X sky130_fd_sc_hd__or2_4
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15587_ _15570_/A _15570_/B _15568_/A vssd1 vssd1 vccd1 vccd1 _15591_/A sky130_fd_sc_hd__o21a_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12795_/X _12798_/X _13130_/A vssd1 vssd1 vccd1 vccd1 _12799_/X sky130_fd_sc_hd__mux2_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17326_ _17326_/A _17326_/B vssd1 vssd1 vccd1 vccd1 _19460_/D sky130_fd_sc_hd__and2_1
XFILLER_30_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14538_ _14596_/A _14538_/B vssd1 vssd1 vccd1 vccd1 _18377_/D sky130_fd_sc_hd__or2_1
XFILLER_159_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17257_ _18113_/Q _17389_/B1 _17453_/A _17256_/B vssd1 vssd1 vccd1 vccd1 _17257_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14469_ _18321_/Q _16540_/A0 _14486_/S vssd1 vssd1 vccd1 vccd1 _18321_/D sky130_fd_sc_hd__mux2_1
X_16208_ _17705_/A0 _18824_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _18824_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17188_ _19414_/Q fanout533/X _17503_/A _17119_/B vssd1 vssd1 vccd1 vccd1 _17189_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_127_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16139_ _18772_/Q _16139_/B vssd1 vssd1 vccd1 vccd1 _16139_/Y sky130_fd_sc_hd__nand2_1
XFILLER_255_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ _11513_/A1 _18318_/Q _17769_/Q _11503_/S0 vssd1 vssd1 vccd1 vccd1 _08961_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08892_ _18112_/Q _11441_/B vssd1 vssd1 vccd1 vccd1 _08892_/X sky130_fd_sc_hd__or2_2
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09513_ _18632_/Q _09883_/B vssd1 vssd1 vccd1 vccd1 _09513_/X sky130_fd_sc_hd__or2_1
XFILLER_271_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09444_ _10315_/S _09442_/X _09443_/X _10996_/B1 vssd1 vssd1 vccd1 vccd1 _09444_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_197_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _10297_/A1 _09370_/X _09371_/X vssd1 vssd1 vccd1 vccd1 _09376_/B sky130_fd_sc_hd__o21ai_1
XFILLER_240_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10150_ _19648_/Q _18937_/Q _10224_/S vssd1 vssd1 vccd1 vccd1 _10150_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput292 _11967_/X vssd1 vssd1 vccd1 vccd1 addr0[7] sky130_fd_sc_hd__buf_4
X_10081_ _15549_/A _11103_/A _09141_/A vssd1 vssd1 vccd1 vccd1 _10081_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13840_ _10905_/S _13810_/A _13839_/X vssd1 vssd1 vccd1 vccd1 _13840_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13771_ _15133_/A _13769_/X _13770_/Y _13869_/B2 vssd1 vssd1 vccd1 vccd1 _13771_/X
+ sky130_fd_sc_hd__a22o_1
X_10983_ _10985_/A _10985_/B vssd1 vssd1 vccd1 vccd1 _10984_/A sky130_fd_sc_hd__and2_1
XFILLER_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15510_ _15487_/A _15487_/B _15485_/Y _15511_/A _15486_/A vssd1 vssd1 vccd1 vccd1
+ _15532_/B sky130_fd_sc_hd__o311a_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12722_ _12721_/X _12720_/X _12821_/A vssd1 vssd1 vccd1 vccd1 _12722_/X sky130_fd_sc_hd__mux2_1
X_16490_ _16490_/A0 _19097_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _19097_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15441_ _15421_/A _15421_/B _15419_/A vssd1 vssd1 vccd1 vccd1 _15445_/A sky130_fd_sc_hd__o21a_2
X_12653_ _10381_/A _12653_/B vssd1 vssd1 vccd1 vccd1 _12653_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_130_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18160_ _19623_/CLK _18160_/D vssd1 vssd1 vccd1 vccd1 _18160_/Q sky130_fd_sc_hd__dfxtp_1
X_11604_ _18470_/Q _18371_/Q _11604_/S vssd1 vssd1 vccd1 vccd1 _11604_/X sky130_fd_sc_hd__mux2_1
X_15372_ _19468_/Q _19402_/Q vssd1 vssd1 vccd1 vccd1 _15373_/B sky130_fd_sc_hd__or2_1
XFILLER_196_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12584_ _12584_/A _12584_/B vssd1 vssd1 vccd1 vccd1 _12584_/Y sky130_fd_sc_hd__nor2_2
X_17111_ _19389_/Q _17115_/B vssd1 vssd1 vccd1 vccd1 _17111_/X sky130_fd_sc_hd__or2_1
X_14323_ _18180_/Q _17707_/A0 _14325_/S vssd1 vssd1 vccd1 vccd1 _18180_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18091_ _18776_/CLK _18091_/D vssd1 vssd1 vccd1 vccd1 _18091_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11535_ _13597_/A _11673_/B _11534_/B _13600_/S vssd1 vssd1 vccd1 vccd1 _11671_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_278_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17042_ _17208_/B _17046_/A2 _17041_/X _17374_/A vssd1 vssd1 vccd1 vccd1 _19357_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14254_ _18125_/Q _14260_/B vssd1 vssd1 vccd1 vccd1 _14254_/X sky130_fd_sc_hd__or2_1
X_11466_ _09129_/S _11464_/X _11465_/X _11466_/B1 vssd1 vssd1 vccd1 vccd1 _11466_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13205_ _17832_/Q _13942_/A2 _13942_/B1 _17864_/Q vssd1 vssd1 vccd1 vccd1 _13205_/X
+ sky130_fd_sc_hd__a22o_1
X_10417_ _18333_/Q _17784_/Q _10426_/S vssd1 vssd1 vccd1 vccd1 _10417_/X sky130_fd_sc_hd__mux2_1
X_11397_ _11397_/A1 _11394_/X _11395_/X _11396_/X vssd1 vssd1 vccd1 vccd1 _11397_/X
+ sky130_fd_sc_hd__a211o_1
X_14185_ _16972_/A _14185_/B vssd1 vssd1 vccd1 vccd1 _18090_/D sky130_fd_sc_hd__and2_1
XFILLER_124_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13136_ _13133_/X _13135_/X _13136_/S vssd1 vssd1 vccd1 vccd1 _13137_/A sky130_fd_sc_hd__mux2_1
X_10348_ _18043_/Q _18011_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _10348_/X sky130_fd_sc_hd__mux2_1
XFILLER_225_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18993_ _19602_/CLK _18993_/D vssd1 vssd1 vccd1 vccd1 _18993_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _19127_/Q _19159_/Q _10281_/S vssd1 vssd1 vccd1 vccd1 _10279_/X sky130_fd_sc_hd__mux2_1
X_17944_ _18627_/CLK _17944_/D vssd1 vssd1 vccd1 vccd1 _17944_/Q sky130_fd_sc_hd__dfxtp_2
X_13067_ _19334_/Q _13246_/A2 _13063_/X _13066_/X _13246_/B1 vssd1 vssd1 vccd1 vccd1
+ _13067_/X sky130_fd_sc_hd__a221o_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1440 _09087_/Y vssd1 vssd1 vccd1 vccd1 _09534_/S sky130_fd_sc_hd__buf_4
X_12018_ _17785_/Q _16553_/A0 _12021_/S vssd1 vssd1 vccd1 vccd1 _17785_/D sky130_fd_sc_hd__mux2_1
X_17875_ _19324_/CLK _17875_/D vssd1 vssd1 vccd1 vccd1 _17875_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1451 _09857_/A1 vssd1 vssd1 vccd1 vccd1 _11156_/C1 sky130_fd_sc_hd__buf_4
Xfanout1462 _10815_/B vssd1 vssd1 vccd1 vccd1 _11598_/S sky130_fd_sc_hd__buf_6
XFILLER_226_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1473 _10511_/S vssd1 vssd1 vccd1 vccd1 _10645_/S sky130_fd_sc_hd__buf_6
XFILLER_238_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1484 fanout1485/X vssd1 vssd1 vccd1 vccd1 _10726_/S sky130_fd_sc_hd__buf_6
XFILLER_266_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19614_ _19614_/CLK _19614_/D vssd1 vssd1 vccd1 vccd1 _19614_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1495 _09428_/B2 vssd1 vssd1 vccd1 vccd1 _10299_/S sky130_fd_sc_hd__buf_6
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16826_ _17810_/Q _14675_/C _16836_/S vssd1 vssd1 vccd1 vccd1 _17118_/B sky130_fd_sc_hd__mux2_2
XFILLER_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16757_ _19272_/Q _16759_/C _16756_/Y vssd1 vssd1 vccd1 vccd1 _19272_/D sky130_fd_sc_hd__a21oi_1
X_19545_ _19546_/CLK _19545_/D vssd1 vssd1 vccd1 vccd1 _19545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13969_ _14268_/A _13969_/B vssd1 vssd1 vccd1 vccd1 _13969_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_81_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15708_ _15789_/A1 _15707_/Y _15789_/B1 vssd1 vssd1 vccd1 vccd1 _15708_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16688_ _19249_/Q _19248_/Q _16688_/C vssd1 vssd1 vccd1 vccd1 _16695_/C sky130_fd_sc_hd__and3_1
X_19476_ _19485_/CLK _19476_/D vssd1 vssd1 vccd1 vccd1 _19476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _15639_/A _15639_/B _15618_/B vssd1 vssd1 vccd1 vccd1 _15640_/B sky130_fd_sc_hd__or3b_1
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18427_ _19575_/CLK _18427_/D vssd1 vssd1 vccd1 vccd1 _18427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09160_ _17930_/Q _08945_/X _09159_/X vssd1 vssd1 vccd1 vccd1 _09160_/X sky130_fd_sc_hd__o21a_4
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18358_ _19636_/CLK _18358_/D vssd1 vssd1 vccd1 vccd1 _18358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17309_ _17307_/Y _17308_/X _17210_/A vssd1 vssd1 vccd1 vccd1 _19453_/D sky130_fd_sc_hd__a21oi_1
X_09091_ _14306_/C _10326_/A vssd1 vssd1 vccd1 vccd1 _09102_/B sky130_fd_sc_hd__nor2_1
X_18289_ _19450_/CLK _18289_/D vssd1 vssd1 vccd1 vccd1 _18289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09993_ _18373_/Q _11692_/A1 _09992_/Y _09043_/A vssd1 vssd1 vccd1 vccd1 _09993_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ _08941_/X _08943_/Y _08940_/X vssd1 vssd1 vccd1 vccd1 _08944_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_269_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08875_ _17914_/Q _17913_/Q _08875_/C _08875_/D vssd1 vssd1 vccd1 vccd1 _08876_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_151_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09427_ _10294_/A1 _19625_/Q _18914_/Q _09428_/B2 vssd1 vssd1 vccd1 vccd1 _09427_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ _11469_/A1 _19139_/Q _09179_/B _19107_/Q _10335_/S vssd1 vssd1 vccd1 vccd1
+ _09358_/X sky130_fd_sc_hd__o221a_1
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09289_ _09284_/X _09288_/X _09958_/C1 vssd1 vssd1 vccd1 vccd1 _09289_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11320_ _11584_/C1 _11317_/X _11318_/X _11319_/X vssd1 vssd1 vccd1 vccd1 _11320_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11251_ _11249_/X _11250_/X _11251_/S vssd1 vssd1 vccd1 vccd1 _11251_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10202_ _18045_/Q _18013_/Q _10206_/S vssd1 vssd1 vccd1 vccd1 _10202_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11182_ _18252_/Q _18827_/Q _18455_/Q _18356_/Q _10717_/S _11199_/S1 vssd1 vssd1
+ vccd1 vccd1 _11183_/B sky130_fd_sc_hd__mux4_1
XFILLER_192_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10133_ _10219_/A1 _18234_/Q _10224_/S _18969_/Q _10225_/S vssd1 vssd1 vccd1 vccd1
+ _10133_/X sky130_fd_sc_hd__o221a_1
XFILLER_267_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15990_ _18710_/Q _16002_/A2 _16004_/B1 _18759_/Q _16004_/C1 vssd1 vssd1 vccd1 vccd1
+ _15990_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14941_ _18495_/Q _14667_/X _14940_/Y _16787_/A vssd1 vssd1 vccd1 vccd1 _18495_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10064_ _12796_/S _12603_/B vssd1 vssd1 vccd1 vccd1 _10065_/B sky130_fd_sc_hd__nand2b_1
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17660_ _17660_/A0 _19587_/Q _17687_/S vssd1 vssd1 vccd1 vccd1 _19587_/D sky130_fd_sc_hd__mux2_1
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14872_ _15003_/A1 _13527_/X _14983_/B1 _18644_/Q _14973_/C1 vssd1 vssd1 vccd1 vccd1
+ _14872_/X sky130_fd_sc_hd__a221o_1
XFILLER_275_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16611_ _16611_/A0 _19214_/Q _16618_/S vssd1 vssd1 vccd1 vccd1 _19214_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13823_ _19549_/Q _13946_/B vssd1 vssd1 vccd1 vccd1 _13823_/X sky130_fd_sc_hd__or2_1
XFILLER_91_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17591_ _17591_/A _17591_/B _17591_/C _17591_/D vssd1 vssd1 vccd1 vccd1 _17591_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_211_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19330_ _19522_/CLK _19330_/D vssd1 vssd1 vccd1 vccd1 _19330_/Q sky130_fd_sc_hd__dfxtp_1
X_16542_ _16542_/A0 _19147_/Q _16548_/S vssd1 vssd1 vccd1 vccd1 _19147_/D sky130_fd_sc_hd__mux2_1
X_13754_ _19321_/Q _13754_/A2 _13747_/X _13753_/X vssd1 vssd1 vccd1 vccd1 _13754_/Y
+ sky130_fd_sc_hd__a211oi_2
X_10966_ _10964_/X _10965_/X _11361_/S vssd1 vssd1 vccd1 vccd1 _10966_/X sky130_fd_sc_hd__mux2_1
XFILLER_245_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19261_ _19261_/CLK _19261_/D vssd1 vssd1 vccd1 vccd1 _19261_/Q sky130_fd_sc_hd__dfxtp_2
X_12705_ _12704_/X _12703_/X _12813_/S vssd1 vssd1 vccd1 vccd1 _12705_/X sky130_fd_sc_hd__mux2_1
X_16473_ _17705_/A0 _19080_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _19080_/D sky130_fd_sc_hd__mux2_1
XFILLER_206_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13685_ _19513_/Q _13947_/A2 _13947_/B1 _13684_/X vssd1 vssd1 vccd1 vccd1 _13685_/X
+ sky130_fd_sc_hd__o211a_1
X_10897_ _10895_/X _10896_/X _11127_/S vssd1 vssd1 vccd1 vccd1 _10897_/X sky130_fd_sc_hd__mux2_1
X_18212_ _19564_/CLK _18212_/D vssd1 vssd1 vccd1 vccd1 _18212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15424_ _17211_/A _15411_/X _15416_/X _15423_/X _15424_/C1 vssd1 vssd1 vccd1 vccd1
+ _15424_/X sky130_fd_sc_hd__a311o_1
XPHY_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19192_ _19647_/CLK _19192_/D vssd1 vssd1 vccd1 vccd1 _19192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12636_ _11676_/A _12593_/Y _13466_/A _12635_/Y vssd1 vssd1 vccd1 vccd1 _13597_/B
+ sky130_fd_sc_hd__a31o_2
XPHY_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18143_ _19203_/CLK _18143_/D vssd1 vssd1 vccd1 vccd1 _18143_/Q sky130_fd_sc_hd__dfxtp_1
X_15355_ _15330_/A _15381_/A3 _15330_/B vssd1 vssd1 vccd1 vccd1 _15484_/A sky130_fd_sc_hd__a21oi_4
XFILLER_184_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12567_ _12768_/B _13167_/B vssd1 vssd1 vccd1 vccd1 _12570_/D sky130_fd_sc_hd__nor2_2
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14306_ _17801_/Q _16392_/B _14306_/C vssd1 vssd1 vccd1 vccd1 _16194_/B sky130_fd_sc_hd__or3_4
X_18074_ _18666_/CLK _18074_/D vssd1 vssd1 vccd1 vccd1 _18074_/Q sky130_fd_sc_hd__dfxtp_1
X_11518_ _11055_/B2 _11517_/X _11452_/B _11518_/B2 vssd1 vssd1 vccd1 vccd1 _15357_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_15286_ _15382_/B2 _15285_/X _15786_/A2 _14224_/A vssd1 vssd1 vccd1 vccd1 _15289_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_12498_ _17823_/Q _13942_/A2 _13942_/B1 _17855_/Q vssd1 vssd1 vccd1 vccd1 _12498_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17025_ _19349_/Q _17045_/B vssd1 vssd1 vccd1 vccd1 _17025_/X sky130_fd_sc_hd__or2_1
X_14237_ _18290_/Q _14261_/A2 _14236_/X _14451_/B vssd1 vssd1 vccd1 vccd1 _18116_/D
+ sky130_fd_sc_hd__o211a_1
X_11449_ _09050_/X _09660_/B _11448_/Y _09030_/X vssd1 vssd1 vccd1 vccd1 _11449_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_171_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14168_ _18695_/Q _18082_/Q _14186_/S vssd1 vssd1 vccd1 vccd1 _14169_/B sky130_fd_sc_hd__mux2_1
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13119_ _12454_/X _13988_/B _13101_/Y vssd1 vssd1 vccd1 vccd1 _13119_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_285_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18976_ _19211_/CLK _18976_/D vssd1 vssd1 vccd1 vccd1 _18976_/Q sky130_fd_sc_hd__dfxtp_1
X_14099_ _17682_/A0 _18039_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _18039_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17927_ _17930_/CLK _17927_/D vssd1 vssd1 vccd1 vccd1 _17927_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1270 _14591_/A2 vssd1 vssd1 vccd1 vccd1 _14575_/A2 sky130_fd_sc_hd__buf_4
Xfanout1281 _15854_/B vssd1 vssd1 vccd1 vccd1 _16016_/A2 sky130_fd_sc_hd__buf_4
XFILLER_67_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17858_ _18691_/CLK _17858_/D vssd1 vssd1 vccd1 vccd1 _17858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1292 _14591_/B1 vssd1 vssd1 vccd1 vccd1 _14589_/B1 sky130_fd_sc_hd__buf_4
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16809_ _19292_/Q _16810_/B vssd1 vssd1 vccd1 vccd1 _16811_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17789_ _19618_/CLK _17789_/D vssd1 vssd1 vccd1 vccd1 _17789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19528_ _19534_/CLK _19528_/D vssd1 vssd1 vccd1 vccd1 _19528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19459_ _19522_/CLK _19459_/D vssd1 vssd1 vccd1 vccd1 _19459_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ _09210_/X _09211_/X _10200_/S vssd1 vssd1 vccd1 vccd1 _09212_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09143_ _09143_/A _12598_/B vssd1 vssd1 vccd1 vccd1 _09145_/A sky130_fd_sc_hd__nor2_2
XFILLER_148_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09074_ _12756_/A _12442_/B vssd1 vssd1 vccd1 vccd1 _12837_/A sky130_fd_sc_hd__nand2_8
XFILLER_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ _09976_/A1 _09969_/X _09968_/X _08967_/S vssd1 vssd1 vccd1 vccd1 _09976_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08927_ _12089_/A _12053_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _08927_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08858_ _08858_/A vssd1 vssd1 vccd1 vccd1 _08858_/Y sky130_fd_sc_hd__inv_2
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10820_ _18460_/Q _18361_/Q _11598_/S vssd1 vssd1 vccd1 vccd1 _10820_/X sky130_fd_sc_hd__mux2_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_98_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19142_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10751_ _18123_/Q _10750_/Y _13739_/A vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__mux2_4
XFILLER_197_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13470_ _12442_/D _13413_/X _13416_/X _12704_/S _13469_/X vssd1 vssd1 vccd1 vccd1
+ _13470_/X sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_27_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19588_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_231_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10682_ _17942_/Q _08948_/B _10681_/X _08947_/B vssd1 vssd1 vccd1 vccd1 _10682_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12421_ _12421_/A _12421_/B vssd1 vssd1 vccd1 vccd1 _12421_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15140_ _19426_/Q _15140_/B vssd1 vssd1 vccd1 vccd1 _15140_/Y sky130_fd_sc_hd__nor2_1
X_12352_ _12379_/A _12352_/B vssd1 vssd1 vccd1 vccd1 _12352_/Y sky130_fd_sc_hd__nand2_1
XFILLER_194_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11303_ _10784_/S _11302_/X _11301_/X _10930_/S vssd1 vssd1 vccd1 vccd1 _11303_/X
+ sky130_fd_sc_hd__a211o_1
X_15071_ _18555_/Q _17682_/A0 _15079_/S vssd1 vssd1 vccd1 vccd1 _18555_/D sky130_fd_sc_hd__mux2_1
X_12283_ _18090_/Q _12305_/A2 _12305_/B1 _18513_/Q vssd1 vssd1 vccd1 vccd1 _12492_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14022_ _17976_/Q _14036_/A vssd1 vssd1 vccd1 vccd1 _14022_/X sky130_fd_sc_hd__or2_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11234_ _11569_/S1 _11233_/X _11232_/X _11248_/S vssd1 vssd1 vccd1 vccd1 _11234_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_162_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18830_ _19637_/CLK _18830_/D vssd1 vssd1 vccd1 vccd1 _18830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11165_ _11480_/C1 _11162_/X _11164_/X vssd1 vssd1 vccd1 vccd1 _11165_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10116_ _18656_/Q _18078_/Q _19097_/Q _19001_/Q _09344_/S _11001_/C1 vssd1 vssd1
+ vccd1 vccd1 _10116_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18761_ _18761_/CLK _18761_/D vssd1 vssd1 vccd1 vccd1 _18761_/Q sky130_fd_sc_hd__dfxtp_2
X_15973_ _18702_/Q _15977_/A2 _15972_/X _16153_/D vssd1 vssd1 vccd1 vccd1 _18702_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_212_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11096_ _11094_/X _11095_/X _11251_/S vssd1 vssd1 vccd1 vccd1 _11096_/X sky130_fd_sc_hd__mux2_1
XFILLER_283_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17712_ _17712_/A0 _19638_/Q _17718_/S vssd1 vssd1 vccd1 vccd1 _19638_/D sky130_fd_sc_hd__mux2_1
X_14924_ _18124_/Q _14893_/S _14852_/X _14923_/X vssd1 vssd1 vccd1 vccd1 _14924_/X
+ sky130_fd_sc_hd__o211a_2
X_10047_ _10045_/X _10046_/X _10719_/S vssd1 vssd1 vccd1 vccd1 _10047_/X sky130_fd_sc_hd__mux2_1
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18692_ _18713_/CLK _18692_/D vssd1 vssd1 vccd1 vccd1 _18692_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_236_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14855_ _14865_/A1 _14853_/X _14865_/B1 vssd1 vssd1 vccd1 vccd1 _14855_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_36_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17643_ _17676_/A0 _19571_/Q _17657_/S vssd1 vssd1 vccd1 vccd1 _19571_/D sky130_fd_sc_hd__mux2_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13806_ _13904_/A _13806_/B vssd1 vssd1 vccd1 vccd1 _13806_/Y sky130_fd_sc_hd__nand2_2
XFILLER_91_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17574_ _19529_/Q _17558_/B _17603_/B1 _17573_/X vssd1 vssd1 vccd1 vccd1 _19529_/D
+ sky130_fd_sc_hd__o211a_1
X_14786_ _14696_/A _18270_/Q _14785_/Y _14846_/B1 vssd1 vssd1 vccd1 vccd1 _14786_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11998_ _17765_/Q _17666_/A0 _12019_/S vssd1 vssd1 vccd1 vccd1 _17765_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19313_ _19363_/CLK _19313_/D vssd1 vssd1 vccd1 vccd1 _19313_/Q sky130_fd_sc_hd__dfxtp_1
X_16525_ _16525_/A _17625_/A vssd1 vssd1 vccd1 vccd1 _16525_/Y sky130_fd_sc_hd__nand2_8
X_13737_ _13802_/C _13737_/B vssd1 vssd1 vccd1 vccd1 _13737_/X sky130_fd_sc_hd__or2_1
X_10949_ _11103_/A _11850_/A vssd1 vssd1 vccd1 vccd1 _10949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19244_ _19280_/CLK _19244_/D vssd1 vssd1 vccd1 vccd1 _19244_/Q sky130_fd_sc_hd__dfxtp_2
X_16456_ _19064_/Q _16621_/A0 _16457_/S vssd1 vssd1 vccd1 vccd1 _19064_/D sky130_fd_sc_hd__mux2_1
X_13668_ _13665_/A _13797_/A0 _13667_/Y _10754_/B vssd1 vssd1 vccd1 vccd1 _13668_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_220_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15407_ _15408_/A _15408_/B vssd1 vssd1 vccd1 vccd1 _15407_/X sky130_fd_sc_hd__or2_2
X_19175_ _19587_/CLK _19175_/D vssd1 vssd1 vccd1 vccd1 _19175_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12619_ _09401_/A _09401_/B _09401_/C vssd1 vssd1 vccd1 vccd1 _13188_/C sky130_fd_sc_hd__o21ba_1
X_16387_ _16553_/A0 _18998_/Q _16390_/S vssd1 vssd1 vccd1 vccd1 _18998_/D sky130_fd_sc_hd__mux2_1
X_13599_ _13611_/B _13961_/A _13598_/X vssd1 vssd1 vccd1 vccd1 _13599_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_247_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18126_ _19450_/CLK _18126_/D vssd1 vssd1 vccd1 vccd1 _18126_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15338_ _15308_/B _15313_/B _15365_/D vssd1 vssd1 vccd1 vccd1 _15340_/A sky130_fd_sc_hd__a21oi_1
XFILLER_172_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18057_ _19140_/CLK _18057_/D vssd1 vssd1 vccd1 vccd1 _18057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15269_ _15267_/X _15268_/Y _15307_/B vssd1 vssd1 vccd1 vccd1 _15274_/B sky130_fd_sc_hd__a21o_1
X_17008_ _17583_/A _17008_/A2 _17007_/X _17342_/A vssd1 vssd1 vccd1 vccd1 _19340_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout507 _17499_/A2 vssd1 vssd1 vccd1 vccd1 _17523_/B sky130_fd_sc_hd__clkbuf_8
X_09830_ _18813_/Q _11224_/B vssd1 vssd1 vccd1 vccd1 _09830_/X sky130_fd_sc_hd__or2_1
Xfanout518 _17241_/B vssd1 vssd1 vccd1 vccd1 _17256_/B sky130_fd_sc_hd__buf_4
Xfanout529 _11770_/B1 vssd1 vssd1 vccd1 vccd1 _11909_/A sky130_fd_sc_hd__buf_2
XFILLER_263_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09761_ _11565_/A1 _18207_/Q _09770_/S _18942_/Q vssd1 vssd1 vccd1 vccd1 _09761_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18959_ _19618_/CLK _18959_/D vssd1 vssd1 vccd1 vccd1 _18959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_273_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09692_ _10180_/A _09670_/X _09691_/X _09686_/Y _09679_/Y vssd1 vssd1 vccd1 vccd1
+ _09692_/X sky130_fd_sc_hd__a32o_2
XFILLER_39_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09126_ _11465_/A1 _18605_/Q _18176_/Q _11455_/S vssd1 vssd1 vccd1 vccd1 _09126_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09057_ _09141_/A _15332_/A _08892_/X vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__o21ai_4
XFILLER_108_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_145_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18778_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_278_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09959_ _12389_/A1 _09949_/X _09950_/X vssd1 vssd1 vccd1 vccd1 _09959_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _19396_/Q _12570_/A _13244_/B1 vssd1 vssd1 vccd1 vccd1 _12970_/X sky130_fd_sc_hd__a21o_1
XFILLER_218_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _11926_/A1 _11939_/A1 _11807_/B _11935_/B1 input226/X vssd1 vssd1 vccd1 vccd1
+ _11921_/X sky130_fd_sc_hd__a32o_4
XFILLER_58_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_401 _09738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_412 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _17699_/A0 _18446_/Q _14660_/S vssd1 vssd1 vccd1 vccd1 _18446_/D sky130_fd_sc_hd__mux2_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_423 _11774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11852_ _11952_/A2 _11850_/X _11851_/X vssd1 vssd1 vccd1 vccd1 _11853_/B sky130_fd_sc_hd__a21oi_4
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_434 _11904_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_445 _14008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_456 _18575_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_467 _18374_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10803_ _11355_/A1 _10802_/X _10801_/X _11338_/S1 vssd1 vssd1 vccd1 vccd1 _10803_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _18394_/Q _14575_/A2 _14575_/B1 input23/X vssd1 vssd1 vccd1 vccd1 _14572_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_478 input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ _11859_/A _11803_/B vssd1 vssd1 vccd1 vccd1 _11783_/Y sky130_fd_sc_hd__nand2_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_489 _18115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16310_ _17708_/A0 _18923_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _18923_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13522_ _19410_/Q _13654_/A2 _13654_/B1 vssd1 vssd1 vccd1 vccd1 _13522_/X sky130_fd_sc_hd__a21o_1
XFILLER_242_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10734_ _19057_/Q _19025_/Q _10744_/S vssd1 vssd1 vccd1 vccd1 _10734_/X sky130_fd_sc_hd__mux2_1
X_17290_ _14252_/A _17199_/A _17508_/A _17289_/B vssd1 vssd1 vccd1 vccd1 _17290_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_213_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16241_ _11376_/B _18856_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _18856_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13453_ _19408_/Q _13654_/A2 _13654_/B1 vssd1 vssd1 vccd1 vccd1 _13453_/X sky130_fd_sc_hd__a21o_1
X_10665_ _10663_/S _10656_/X _10657_/X vssd1 vssd1 vccd1 vccd1 _10665_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12404_ _12471_/A0 _12430_/A _12403_/Y _14001_/C1 vssd1 vssd1 vccd1 vccd1 _17909_/D
+ sky130_fd_sc_hd__o211a_1
X_16172_ _16602_/A0 _18789_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _18789_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13384_ _13791_/A _13382_/Y _13383_/X _13402_/B _13622_/A vssd1 vssd1 vccd1 vccd1
+ _13384_/X sky130_fd_sc_hd__a32o_1
XFILLER_154_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ _11602_/C1 _10589_/X _11608_/C1 vssd1 vssd1 vccd1 vccd1 _10596_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_166_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15123_ _17124_/A _15123_/B _15118_/Y vssd1 vssd1 vccd1 vccd1 _15123_/X sky130_fd_sc_hd__or3b_1
X_12335_ _17796_/Q _08905_/X _08939_/A _08942_/Y _12334_/Y vssd1 vssd1 vccd1 vccd1
+ _12335_/X sky130_fd_sc_hd__a41o_2
XFILLER_127_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15054_ _18538_/Q _16532_/A0 _15076_/S vssd1 vssd1 vccd1 vccd1 _18538_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12266_ _17891_/Q _17890_/Q vssd1 vssd1 vccd1 vccd1 _12267_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14005_ _17967_/Q _14036_/A _14004_/Y _14037_/C1 vssd1 vssd1 vccd1 vccd1 _17967_/D
+ sky130_fd_sc_hd__o211a_1
X_11217_ _11217_/A _11217_/B _11217_/C vssd1 vssd1 vccd1 vccd1 _11217_/X sky130_fd_sc_hd__and3_1
XFILLER_268_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12197_ _17863_/Q _12200_/C _12203_/A vssd1 vssd1 vccd1 vccd1 _12197_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_269_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18813_ _19195_/CLK _18813_/D vssd1 vssd1 vccd1 vccd1 _18813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11148_ _11567_/S _11147_/X _11146_/X _09845_/S vssd1 vssd1 vccd1 vccd1 _11148_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_268_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18744_ _18746_/CLK _18744_/D vssd1 vssd1 vccd1 vccd1 _18744_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_283_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15956_ _15854_/A _15970_/A2 _15976_/B1 _18742_/Q _15976_/C1 vssd1 vssd1 vccd1 vccd1
+ _15956_/X sky130_fd_sc_hd__a221o_1
X_11079_ _11305_/A1 _19571_/Q _11309_/S _19603_/Q _11311_/C1 vssd1 vssd1 vccd1 vccd1
+ _11079_/X sky130_fd_sc_hd__o221a_1
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput170 dout1[9] vssd1 vssd1 vccd1 vccd1 input170/X sky130_fd_sc_hd__clkbuf_2
XFILLER_271_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput181 irq[4] vssd1 vssd1 vccd1 vccd1 _15084_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput192 localMemory_wb_adr_i[11] vssd1 vssd1 vccd1 vccd1 input192/X sky130_fd_sc_hd__clkbuf_2
X_14907_ _14907_/A vssd1 vssd1 vccd1 vccd1 _14907_/Y sky130_fd_sc_hd__clkinv_4
X_18675_ _18683_/CLK _18675_/D vssd1 vssd1 vccd1 vccd1 _18675_/Q sky130_fd_sc_hd__dfxtp_1
X_15887_ _15887_/A _15905_/B _15923_/C vssd1 vssd1 vccd1 vccd1 _15887_/X sky130_fd_sc_hd__and3_1
XFILLER_236_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17626_ _17659_/A0 _19554_/Q _17648_/S vssd1 vssd1 vccd1 vccd1 _19554_/D sky130_fd_sc_hd__mux2_1
X_14838_ _18485_/Q _15001_/A2 _14837_/Y _16808_/A vssd1 vssd1 vccd1 vccd1 _18485_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14769_ _14973_/A1 _13180_/Y _14973_/B1 _18634_/Q _14741_/B vssd1 vssd1 vccd1 vccd1
+ _14769_/X sky130_fd_sc_hd__a221o_2
X_17557_ _17559_/B _17583_/B vssd1 vssd1 vccd1 vccd1 _17557_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16508_ _17674_/A0 _19114_/Q _16515_/S vssd1 vssd1 vccd1 vccd1 _19114_/D sky130_fd_sc_hd__mux2_1
X_17488_ _17488_/A _17493_/B vssd1 vssd1 vccd1 vccd1 _17488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19227_ _19229_/CLK _19227_/D vssd1 vssd1 vccd1 vccd1 _19227_/Q sky130_fd_sc_hd__dfxtp_4
X_16439_ _19047_/Q _11452_/B _16454_/S vssd1 vssd1 vccd1 vccd1 _19047_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19158_ _19596_/CLK _19158_/D vssd1 vssd1 vccd1 vccd1 _19158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18109_ _19448_/CLK _18109_/D vssd1 vssd1 vccd1 vccd1 _18109_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_258_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19089_ _19211_/CLK _19089_/D vssd1 vssd1 vccd1 vccd1 _19089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09813_ _11210_/A1 _09743_/B _09812_/X _11055_/B2 vssd1 vssd1 vccd1 vccd1 _15151_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09744_ _18846_/Q _18878_/Q _09770_/S vssd1 vssd1 vccd1 vccd1 _09744_/X sky130_fd_sc_hd__mux2_1
XFILLER_246_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09675_ _11172_/A1 _19558_/Q _09688_/S _19590_/Q vssd1 vssd1 vccd1 vccd1 _09675_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10450_ _13775_/A vssd1 vssd1 vccd1 vccd1 _10450_/Y sky130_fd_sc_hd__inv_2
X_09109_ _12468_/B _18144_/Q _18790_/Q _09539_/S _09683_/A vssd1 vssd1 vccd1 vccd1
+ _09109_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10381_ _10381_/A _12653_/B vssd1 vssd1 vccd1 vccd1 _11550_/B sky130_fd_sc_hd__and2_4
XFILLER_151_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12120_ _17833_/Q _17834_/Q _12120_/C vssd1 vssd1 vccd1 vccd1 _12122_/B sky130_fd_sc_hd__and3_1
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12051_ _12051_/A _12051_/B vssd1 vssd1 vccd1 vccd1 _12051_/X sky130_fd_sc_hd__or2_1
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1803 _14427_/B vssd1 vssd1 vccd1 vccd1 _16052_/A sky130_fd_sc_hd__buf_4
X_11002_ _11389_/A1 _17776_/Q _11386_/S _18325_/Q _11002_/C1 vssd1 vssd1 vccd1 vccd1
+ _11002_/X sky130_fd_sc_hd__o221a_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1814 _17354_/A vssd1 vssd1 vccd1 vccd1 _17356_/A sky130_fd_sc_hd__buf_4
XFILLER_105_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1825 _17350_/A vssd1 vssd1 vccd1 vccd1 _17352_/A sky130_fd_sc_hd__buf_4
XFILLER_42_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1836 _14417_/A vssd1 vssd1 vccd1 vccd1 _13981_/C1 sky130_fd_sc_hd__buf_4
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1847 _17342_/A vssd1 vssd1 vccd1 vccd1 _17559_/A sky130_fd_sc_hd__buf_4
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1858 fanout1863/X vssd1 vssd1 vccd1 vccd1 _14001_/C1 sky130_fd_sc_hd__buf_4
Xfanout860 _16615_/A0 vssd1 vssd1 vccd1 vccd1 _17715_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1869 fanout1870/X vssd1 vssd1 vccd1 vccd1 _16812_/B1 sky130_fd_sc_hd__clkbuf_4
X_15810_ _18602_/Q _16203_/A0 _15829_/S vssd1 vssd1 vccd1 vccd1 _18602_/D sky130_fd_sc_hd__mux2_1
Xfanout871 _10239_/B vssd1 vssd1 vccd1 vccd1 _16488_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_77_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16790_ _19284_/Q _16791_/C _19285_/Q vssd1 vssd1 vccd1 vccd1 _16792_/B sky130_fd_sc_hd__a21oi_1
XFILLER_237_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout882 _12818_/S vssd1 vssd1 vccd1 vccd1 _12823_/A sky130_fd_sc_hd__buf_4
Xfanout893 _13039_/S vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__buf_4
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15741_ _18590_/Q _15800_/A2 _15733_/Y _15740_/X _14449_/B vssd1 vssd1 vccd1 vccd1
+ _18590_/D sky130_fd_sc_hd__o221a_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _13315_/S _12952_/Y _13197_/B1 vssd1 vssd1 vccd1 vccd1 _12953_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _11909_/A _11904_/B vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_42_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18902_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15672_ _15672_/A _15672_/B vssd1 vssd1 vccd1 vccd1 _15673_/B sky130_fd_sc_hd__xnor2_1
X_18460_ _19216_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12884_ _12722_/X _12735_/Y _12942_/S vssd1 vssd1 vccd1 vccd1 _12885_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_220 _18640_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_231 _18390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_242 _18380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14623_ _17682_/A0 _18430_/Q _14631_/S vssd1 vssd1 vccd1 vccd1 _18430_/D sky130_fd_sc_hd__mux2_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _18566_/Q _17461_/A2 _17426_/B1 vssd1 vssd1 vccd1 vccd1 _17411_/X sky130_fd_sc_hd__o21a_1
XFILLER_260_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11835_ _14141_/B _11833_/A _11834_/Y _11810_/A vssd1 vssd1 vccd1 vccd1 _11836_/B
+ sky130_fd_sc_hd__o211a_4
XANTENNA_253 _15087_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18391_ _19465_/CLK _18391_/D vssd1 vssd1 vccd1 vccd1 _18391_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 input224/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_275 input240/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 _11890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17342_/A _17342_/B vssd1 vssd1 vccd1 vccd1 _19468_/D sky130_fd_sc_hd__and2_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_297 _18734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14586_/A _14554_/B vssd1 vssd1 vccd1 vccd1 _18385_/D sky130_fd_sc_hd__or2_1
XFILLER_187_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _18584_/Q _14349_/B _11769_/B1 _11686_/A vssd1 vssd1 vccd1 vccd1 _11766_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _14008_/B vssd1 vssd1 vccd1 vccd1 _13505_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10717_ _18329_/Q _17780_/Q _10717_/S vssd1 vssd1 vccd1 vccd1 _10717_/X sky130_fd_sc_hd__mux2_1
X_17273_ _17271_/Y _17272_/X _14423_/B vssd1 vssd1 vccd1 vccd1 _19441_/D sky130_fd_sc_hd__a21oi_1
X_14485_ _18337_/Q _17722_/A0 _14485_/S vssd1 vssd1 vccd1 vccd1 _18337_/D sky130_fd_sc_hd__mux2_1
X_11697_ _11687_/Y _11692_/X _11694_/Y _11695_/X _12461_/A vssd1 vssd1 vccd1 vccd1
+ _11697_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_158_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16224_ _17721_/A0 _18840_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _18840_/D sky130_fd_sc_hd__mux2_1
X_19012_ _19208_/CLK _19012_/D vssd1 vssd1 vccd1 vccd1 _19012_/Q sky130_fd_sc_hd__dfxtp_1
X_13436_ _14004_/B vssd1 vssd1 vccd1 vccd1 _13436_/Y sky130_fd_sc_hd__inv_2
X_10648_ _19122_/Q _19154_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _10648_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16155_ _18275_/D _16156_/B vssd1 vssd1 vccd1 vccd1 _16155_/X sky130_fd_sc_hd__and2_1
X_13367_ _17901_/Q _12448_/C _13365_/Y _13366_/X _12762_/B vssd1 vssd1 vccd1 vccd1
+ _13367_/X sky130_fd_sc_hd__a221o_4
X_10579_ _10881_/S1 _10568_/X _10578_/X _11621_/C1 vssd1 vssd1 vccd1 vccd1 _10579_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _09095_/A _12318_/Y _15285_/A3 _08853_/Y vssd1 vssd1 vccd1 vccd1 _15108_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_142_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12318_ _12318_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _12318_/Y sky130_fd_sc_hd__nor2_2
X_16086_ _16096_/A1 _16085_/Y _17725_/C1 vssd1 vssd1 vccd1 vccd1 _18745_/D sky130_fd_sc_hd__a21oi_1
XFILLER_154_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13298_ _19534_/Q _19502_/Q _13372_/S vssd1 vssd1 vccd1 vccd1 _13298_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ _18526_/Q _12269_/C _15037_/S vssd1 vssd1 vccd1 vccd1 _18526_/D sky130_fd_sc_hd__mux2_1
X_12249_ _12249_/A _12249_/B _12253_/C vssd1 vssd1 vccd1 vccd1 _17882_/D sky130_fd_sc_hd__nor3_1
XFILLER_69_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16988_ _17563_/A _17044_/A2 _16987_/X _17378_/A vssd1 vssd1 vccd1 vccd1 _19330_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18727_ _18734_/CLK _18727_/D vssd1 vssd1 vccd1 vccd1 _18727_/Q sky130_fd_sc_hd__dfxtp_1
X_15939_ _18688_/Q _15948_/A2 _15948_/B1 _15938_/X _15948_/C1 vssd1 vssd1 vccd1 vccd1
+ _15939_/X sky130_fd_sc_hd__a221o_1
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09460_ _09690_/A _09454_/X _09459_/X _08843_/A vssd1 vssd1 vccd1 vccd1 _09460_/X
+ sky130_fd_sc_hd__o211a_1
X_18658_ _18660_/CLK _18658_/D vssd1 vssd1 vccd1 vccd1 _18658_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17609_ _19384_/Q _15088_/B input185/X _17592_/X _17623_/B1 vssd1 vssd1 vccd1 vccd1
+ _17609_/X sky130_fd_sc_hd__a41o_1
XFILLER_251_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09391_ _09389_/X _09390_/X _10225_/S vssd1 vssd1 vccd1 vccd1 _09391_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18589_ _19482_/CLK _18589_/D vssd1 vssd1 vccd1 vccd1 _18589_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_212_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput430 _18499_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[28] sky130_fd_sc_hd__buf_4
Xoutput441 _18480_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[9] sky130_fd_sc_hd__buf_4
XFILLER_105_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput452 _18112_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[11] sky130_fd_sc_hd__buf_4
XFILLER_105_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput463 _18122_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[21] sky130_fd_sc_hd__buf_4
Xoutput474 _18132_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[31] sky130_fd_sc_hd__buf_4
Xoutput485 _11955_/X vssd1 vssd1 vccd1 vccd1 wmask0[1] sky130_fd_sc_hd__buf_4
XFILLER_160_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09727_ _09718_/S _09720_/X _09719_/X _09429_/S vssd1 vssd1 vccd1 vccd1 _09727_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09658_ _09908_/A1 _09236_/A _09657_/X _09908_/B1 _18393_/Q vssd1 vssd1 vccd1 vccd1
+ _09658_/X sky130_fd_sc_hd__o32a_1
XFILLER_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09589_ _19623_/Q _18912_/Q _10370_/S vssd1 vssd1 vccd1 vccd1 _09589_/X sky130_fd_sc_hd__mux2_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11611_/S _11613_/X _11612_/X _11127_/S vssd1 vssd1 vccd1 vccd1 _11620_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11551_ _13794_/A _11639_/B _13812_/A _11549_/X vssd1 vssd1 vccd1 vccd1 _11637_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10502_ _10643_/S _10500_/X _10501_/X _10653_/C1 vssd1 vssd1 vccd1 vccd1 _10502_/X
+ sky130_fd_sc_hd__a211o_1
X_14270_ _16392_/B _16392_/C _17800_/Q vssd1 vssd1 vccd1 vccd1 _16260_/B sky130_fd_sc_hd__and3b_2
X_11482_ _18145_/Q _11482_/A2 _11481_/X _12488_/B vssd1 vssd1 vccd1 vccd1 _11482_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_137_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_160_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19543_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13221_ _15330_/A _13203_/A _13220_/X _13199_/X _13237_/B1 vssd1 vssd1 vccd1 vccd1
+ _13221_/Y sky130_fd_sc_hd__o2111ai_2
X_10433_ _11596_/A1 _19221_/Q _19189_/Q _10815_/B _08899_/A vssd1 vssd1 vccd1 vccd1
+ _10433_/X sky130_fd_sc_hd__a221o_1
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13152_ _13152_/A vssd1 vssd1 vccd1 vccd1 _13152_/Y sky130_fd_sc_hd__inv_2
X_10364_ _18902_/Q _10364_/B vssd1 vssd1 vccd1 vccd1 _10364_/X sky130_fd_sc_hd__or2_1
XFILLER_163_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _17828_/Q _12106_/C vssd1 vssd1 vccd1 vccd1 _12104_/B sky130_fd_sc_hd__and2_1
XFILLER_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17960_ _17982_/CLK _17960_/D vssd1 vssd1 vccd1 vccd1 _17960_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13083_ _13083_/A _13083_/B _13083_/C vssd1 vssd1 vccd1 vccd1 _13084_/B sky130_fd_sc_hd__nand3_1
X_10295_ _10292_/X _10293_/X _10294_/X _10297_/A1 _10301_/S vssd1 vssd1 vccd1 vccd1
+ _10295_/X sky130_fd_sc_hd__a221o_1
XFILLER_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16911_ _19312_/Q _17169_/B _16947_/S vssd1 vssd1 vccd1 vccd1 _16912_/B sky130_fd_sc_hd__mux2_1
Xfanout1600 _08893_/Y vssd1 vssd1 vccd1 vccd1 _11516_/B1 sky130_fd_sc_hd__clkbuf_16
X_12034_ _17892_/Q _12052_/A2 _12033_/X _12383_/C1 vssd1 vssd1 vccd1 vccd1 _17794_/D
+ sky130_fd_sc_hd__o211a_1
Xfanout1611 _16137_/B vssd1 vssd1 vccd1 vccd1 _16141_/B sky130_fd_sc_hd__buf_4
Xfanout1622 _09007_/Y vssd1 vssd1 vccd1 vccd1 _12409_/A2 sky130_fd_sc_hd__buf_4
X_17891_ _17901_/CLK _17891_/D vssd1 vssd1 vccd1 vccd1 _17891_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1633 _15082_/A vssd1 vssd1 vccd1 vccd1 _12023_/A sky130_fd_sc_hd__buf_12
XFILLER_120_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1644 _10817_/A1 vssd1 vssd1 vccd1 vccd1 _11594_/A1 sky130_fd_sc_hd__clkbuf_8
X_19630_ _19630_/CLK _19630_/D vssd1 vssd1 vccd1 vccd1 _19630_/Q sky130_fd_sc_hd__dfxtp_1
X_16842_ _17316_/A vssd1 vssd1 vccd1 vccd1 _16843_/D sky130_fd_sc_hd__inv_2
Xfanout1655 _09873_/A1 vssd1 vssd1 vccd1 vccd1 _10282_/A1 sky130_fd_sc_hd__buf_6
Xfanout1666 _10030_/C1 vssd1 vssd1 vccd1 vccd1 _12766_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_66_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1677 _11584_/A1 vssd1 vssd1 vccd1 vccd1 _10850_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_281_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1688 _10262_/A1 vssd1 vssd1 vccd1 vccd1 _10263_/A1 sky130_fd_sc_hd__buf_6
Xfanout690 _12558_/Y vssd1 vssd1 vccd1 vccd1 _13244_/B1 sky130_fd_sc_hd__buf_6
XFILLER_19_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1699 _09095_/A vssd1 vssd1 vccd1 vccd1 _11584_/C1 sky130_fd_sc_hd__buf_8
XFILLER_253_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19561_ _19614_/CLK _19561_/D vssd1 vssd1 vccd1 vccd1 _19561_/Q sky130_fd_sc_hd__dfxtp_1
X_16773_ _19278_/Q _16775_/C _16772_/Y vssd1 vssd1 vccd1 vccd1 _19278_/D sky130_fd_sc_hd__a21oi_1
X_13985_ _14033_/A1 _13024_/X _13984_/X _14417_/A vssd1 vssd1 vccd1 vccd1 _17957_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18512_ _19321_/CLK _18512_/D vssd1 vssd1 vccd1 vccd1 _18512_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_206_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12936_ _12934_/Y _12935_/X _12936_/S vssd1 vssd1 vccd1 vccd1 _13263_/B sky130_fd_sc_hd__mux2_1
X_15724_ _15724_/A vssd1 vssd1 vccd1 vccd1 _15728_/A sky130_fd_sc_hd__inv_2
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19492_ _19492_/CLK _19492_/D vssd1 vssd1 vccd1 vccd1 _19492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18443_ _19622_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15655_ _15717_/B2 _15654_/X _15782_/B1 vssd1 vssd1 vccd1 vccd1 _15655_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _13438_/A _12847_/X _13956_/B1 vssd1 vssd1 vccd1 vccd1 _12867_/X sky130_fd_sc_hd__a21o_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _16532_/A0 _18413_/Q _14628_/S vssd1 vssd1 vccd1 vccd1 _18413_/D sky130_fd_sc_hd__mux2_1
X_11818_ _11818_/A _11818_/B _11818_/C vssd1 vssd1 vccd1 vccd1 _11818_/X sky130_fd_sc_hd__and3_1
X_15586_ _19445_/Q _15793_/A2 _17199_/A _15585_/X vssd1 vssd1 vccd1 vccd1 _15586_/X
+ sky130_fd_sc_hd__o211a_1
X_18374_ _19465_/CLK _18374_/D vssd1 vssd1 vccd1 vccd1 _18374_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_199_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12798_ _12796_/X _12797_/X _12942_/S vssd1 vssd1 vccd1 vccd1 _12798_/X sky130_fd_sc_hd__mux2_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _19460_/Q _17567_/A _17345_/S vssd1 vssd1 vccd1 vccd1 _17326_/B sky130_fd_sc_hd__mux2_1
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14537_ _18377_/Q _14559_/A2 _14559_/B1 input36/X vssd1 vssd1 vccd1 vccd1 _14538_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11749_ _18570_/Q _14522_/A2 _11818_/B _13147_/A vssd1 vssd1 vccd1 vccd1 _11749_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14468_ _18320_/Q _17672_/A0 _14485_/S vssd1 vssd1 vccd1 vccd1 _18320_/D sky130_fd_sc_hd__mux2_1
X_17256_ _19436_/Q _17256_/B vssd1 vssd1 vccd1 vccd1 _17256_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16207_ _17704_/A0 _18823_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _18823_/D sky130_fd_sc_hd__mux2_1
X_13419_ _12835_/A _13413_/X _13416_/X _12442_/D _13418_/X vssd1 vssd1 vccd1 vccd1
+ _13419_/X sky130_fd_sc_hd__o221a_1
X_17187_ _17202_/A _17187_/B vssd1 vssd1 vccd1 vccd1 _17503_/A sky130_fd_sc_hd__nand2_2
X_14399_ _16606_/A0 _18250_/Q _14416_/S vssd1 vssd1 vccd1 vccd1 _18250_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16138_ _16078_/X _16137_/Y _16142_/B1 vssd1 vssd1 vccd1 vccd1 _18771_/D sky130_fd_sc_hd__a21oi_1
XFILLER_6_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08960_ _11513_/A1 _19597_/Q _19565_/Q _11503_/S0 vssd1 vssd1 vccd1 vccd1 _08960_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16069_ _16069_/A _16069_/B vssd1 vssd1 vccd1 vccd1 _16075_/C sky130_fd_sc_hd__or2_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08891_ _17894_/Q _17893_/Q _09070_/D _12439_/A vssd1 vssd1 vccd1 vccd1 _13807_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_284_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09512_ _18022_/Q _17990_/Q _09724_/S vssd1 vssd1 vccd1 vccd1 _09512_/X sky130_fd_sc_hd__mux2_1
XFILLER_271_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09443_ _10263_/A1 _19138_/Q _09671_/S _19106_/Q _10264_/S vssd1 vssd1 vccd1 vccd1
+ _09443_/X sky130_fd_sc_hd__o221a_1
XFILLER_64_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09374_ _09372_/X _09373_/X _09374_/S vssd1 vssd1 vccd1 vccd1 _09374_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput293 _11968_/X vssd1 vssd1 vccd1 vccd1 addr0[8] sky130_fd_sc_hd__buf_4
X_10080_ _13261_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _13258_/A sky130_fd_sc_hd__xnor2_4
XFILLER_248_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13770_ _18126_/Q _13802_/C vssd1 vssd1 vccd1 vccd1 _13770_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_261_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10982_ _10985_/B vssd1 vssd1 vccd1 vccd1 _10982_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12721_ _10985_/B _11522_/B _12721_/S vssd1 vssd1 vccd1 vccd1 _12721_/X sky130_fd_sc_hd__mux2_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15440_ _19471_/Q _15498_/S vssd1 vssd1 vccd1 vccd1 _15440_/Y sky130_fd_sc_hd__nor2_1
X_12652_ _11639_/A _12651_/X _12648_/X vssd1 vssd1 vccd1 vccd1 _12652_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ _10036_/S _11593_/X _11594_/X vssd1 vssd1 vccd1 vccd1 _11603_/X sky130_fd_sc_hd__o21a_1
X_15371_ _19468_/Q _19402_/Q vssd1 vssd1 vccd1 vccd1 _15373_/A sky130_fd_sc_hd__nand2_2
X_12583_ _13165_/C _12584_/B vssd1 vssd1 vccd1 vccd1 _12583_/Y sky130_fd_sc_hd__nor2_8
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14322_ _18179_/Q _16606_/A0 _14339_/S vssd1 vssd1 vccd1 vccd1 _18179_/D sky130_fd_sc_hd__mux2_1
X_17110_ _17205_/B _17116_/A2 _17109_/X _17368_/A vssd1 vssd1 vccd1 vccd1 _19388_/D
+ sky130_fd_sc_hd__o211a_1
X_18090_ _18776_/CLK _18090_/D vssd1 vssd1 vccd1 vccd1 _18090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11534_ _11673_/B _11534_/B vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__nand2_2
XFILLER_129_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17041_ _19357_/Q _17041_/B vssd1 vssd1 vccd1 vccd1 _17041_/X sky130_fd_sc_hd__or2_1
XFILLER_239_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14253_ _18298_/Q _14252_/B _14252_/Y _17376_/A vssd1 vssd1 vccd1 vccd1 _18124_/D
+ sky130_fd_sc_hd__o211a_1
X_11465_ _11465_/A1 _17770_/Q _11462_/S _18319_/Q _10408_/S vssd1 vssd1 vccd1 vccd1
+ _11465_/X sky130_fd_sc_hd__o221a_1
XFILLER_183_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13204_ _15284_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__and2_1
X_10416_ _17914_/Q _11490_/B _11489_/B1 _10415_/Y vssd1 vssd1 vccd1 vccd1 _10453_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14184_ _18703_/Q _18090_/Q _14186_/S vssd1 vssd1 vccd1 vccd1 _14185_/B sky130_fd_sc_hd__mux2_1
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11396_ _11481_/A _11404_/A1 _19208_/Q _11406_/B2 vssd1 vssd1 vccd1 vccd1 _11396_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13135_ _12750_/X _13414_/B _13135_/S vssd1 vssd1 vccd1 vccd1 _13135_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10347_ _10354_/A1 _19581_/Q _10348_/S _19613_/Q _10205_/S vssd1 vssd1 vccd1 vccd1
+ _10347_/X sky130_fd_sc_hd__o221a_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ _19226_/CLK _18992_/D vssd1 vssd1 vccd1 vccd1 _18992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17943_ _17975_/CLK _17943_/D vssd1 vssd1 vccd1 vccd1 _17943_/Q sky130_fd_sc_hd__dfxtp_2
X_13066_ _19398_/Q _12570_/A _13064_/X _13065_/X _13244_/B1 vssd1 vssd1 vccd1 vccd1
+ _13066_/X sky130_fd_sc_hd__a221o_1
XFILLER_140_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10278_ _18654_/Q _18076_/Q _10281_/S vssd1 vssd1 vccd1 vccd1 _10278_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12017_ _17784_/Q _17685_/A0 _12021_/S vssd1 vssd1 vccd1 vccd1 _17784_/D sky130_fd_sc_hd__mux2_1
Xfanout1430 _10326_/A vssd1 vssd1 vccd1 vccd1 _10623_/A sky130_fd_sc_hd__buf_4
Xfanout1441 _09935_/A vssd1 vssd1 vccd1 vccd1 _10264_/S sky130_fd_sc_hd__buf_8
XFILLER_66_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17874_ _19324_/CLK _17874_/D vssd1 vssd1 vccd1 vccd1 _17874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1452 _09086_/Y vssd1 vssd1 vccd1 vccd1 _09857_/A1 sky130_fd_sc_hd__buf_4
XFILLER_266_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1463 _11360_/B2 vssd1 vssd1 vccd1 vccd1 _10815_/B sky130_fd_sc_hd__buf_6
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19613_ _19613_/CLK _19613_/D vssd1 vssd1 vccd1 vccd1 _19613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1474 _10511_/S vssd1 vssd1 vccd1 vccd1 _10650_/S sky130_fd_sc_hd__buf_4
XFILLER_238_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16825_ _16836_/S _17816_/Q _12478_/Y vssd1 vssd1 vccd1 vccd1 _17051_/A sky130_fd_sc_hd__o21ba_4
XFILLER_94_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1485 fanout1525/X vssd1 vssd1 vccd1 vccd1 fanout1485/X sky130_fd_sc_hd__buf_4
XFILLER_285_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1496 _10290_/S vssd1 vssd1 vccd1 vccd1 _09428_/B2 sky130_fd_sc_hd__buf_6
XFILLER_19_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19544_ _19553_/CLK _19544_/D vssd1 vssd1 vccd1 vccd1 _19544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16756_ _19272_/Q _16759_/C _16764_/B1 vssd1 vssd1 vccd1 vccd1 _16756_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_235_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13968_ _13968_/A1 _13957_/X _13967_/X _13968_/B2 vssd1 vssd1 vccd1 vccd1 _13968_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15707_ _15707_/A _15707_/B vssd1 vssd1 vccd1 vccd1 _15707_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12919_ _17858_/Q _12919_/A2 _12908_/X _13303_/B2 _12918_/X vssd1 vssd1 vccd1 vccd1
+ _12919_/X sky130_fd_sc_hd__a221o_1
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19475_ _19519_/CLK _19475_/D vssd1 vssd1 vccd1 vccd1 _19475_/Q sky130_fd_sc_hd__dfxtp_1
X_16687_ _19248_/Q _16688_/C _16686_/Y vssd1 vssd1 vccd1 vccd1 _19248_/D sky130_fd_sc_hd__o21a_1
X_13899_ _13899_/A _13899_/B vssd1 vssd1 vccd1 vccd1 _13899_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18426_ _18613_/CLK _18426_/D vssd1 vssd1 vccd1 vccd1 _18426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15638_ _15638_/A _15638_/B _15638_/C _15638_/D vssd1 vssd1 vccd1 vccd1 _15638_/X
+ sky130_fd_sc_hd__or4_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18357_ _19637_/CLK _18357_/D vssd1 vssd1 vccd1 vccd1 _18357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15569_ _15540_/Y _15544_/B _15542_/B vssd1 vssd1 vccd1 vccd1 _15570_/B sky130_fd_sc_hd__o21a_1
XFILLER_221_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17308_ _18130_/Q _15782_/A1 _17208_/Y _17307_/B vssd1 vssd1 vccd1 vccd1 _17308_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09090_ _14488_/C _09107_/D vssd1 vssd1 vccd1 vccd1 _09102_/A sky130_fd_sc_hd__nor2_1
X_18288_ _19450_/CLK _18288_/D vssd1 vssd1 vccd1 vccd1 _18288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17239_ _18107_/Q _17382_/A _17423_/A _17241_/B vssd1 vssd1 vccd1 vccd1 _17239_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_163_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09992_ _09992_/A _09992_/B vssd1 vssd1 vccd1 vccd1 _09992_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08943_ _17793_/Q _08927_/Y _08942_/Y _17796_/Q vssd1 vssd1 vccd1 vccd1 _08943_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_142_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08874_ _11252_/S _09777_/A _17906_/Q _08874_/D vssd1 vssd1 vccd1 vccd1 _08875_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09426_ _09718_/S _09426_/B vssd1 vssd1 vccd1 vccd1 _09426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09357_ _11469_/A1 _18212_/Q _09179_/B _18947_/Q _11001_/C1 vssd1 vssd1 vccd1 vccd1
+ _09357_/X sky130_fd_sc_hd__o221a_1
XFILLER_212_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09288_ _09967_/S _09287_/X _09286_/X _10301_/S vssd1 vssd1 vccd1 vccd1 _09288_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ _11250_/A1 _18148_/Q _18794_/Q _11249_/S vssd1 vssd1 vccd1 vccd1 _11250_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10201_ _10354_/A1 _19583_/Q _10199_/S _19615_/Q _10205_/S vssd1 vssd1 vccd1 vccd1
+ _10201_/X sky130_fd_sc_hd__o221a_1
XFILLER_162_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11181_ _10513_/S _11337_/B _11181_/B1 _11180_/Y vssd1 vssd1 vccd1 vccd1 _11214_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10132_ _19097_/Q _19001_/Q _10224_/S vssd1 vssd1 vccd1 vccd1 _10132_/X sky130_fd_sc_hd__mux2_1
XFILLER_267_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14940_ _14936_/Y _14939_/X _15010_/B1 vssd1 vssd1 vccd1 vccd1 _14940_/Y sky130_fd_sc_hd__a21oi_4
X_10063_ _12796_/S _12603_/B vssd1 vssd1 vccd1 vccd1 _11651_/B sky130_fd_sc_hd__and2b_1
XFILLER_134_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ _17808_/Q _14911_/B vssd1 vssd1 vccd1 vccd1 _14871_/X sky130_fd_sc_hd__or2_1
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16610_ _16610_/A0 _19213_/Q _16622_/S vssd1 vssd1 vccd1 vccd1 _19213_/D sky130_fd_sc_hd__mux2_1
XFILLER_217_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13822_ _17882_/Q _13847_/A2 _13820_/X _13920_/B2 vssd1 vssd1 vccd1 vccd1 _13822_/X
+ sky130_fd_sc_hd__a22o_1
X_17590_ _19537_/Q _17622_/A2 _17623_/B1 _17589_/X vssd1 vssd1 vccd1 vccd1 _19537_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13753_ _19385_/Q _13884_/A2 _13751_/X _13752_/X _13884_/C1 vssd1 vssd1 vccd1 vccd1
+ _13753_/X sky130_fd_sc_hd__o221a_4
X_16541_ _17674_/A0 _19146_/Q _16548_/S vssd1 vssd1 vccd1 vccd1 _19146_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10965_ _11596_/A1 _18152_/Q _18798_/Q _11340_/B2 vssd1 vssd1 vccd1 vccd1 _10965_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12704_ _09896_/Y _12657_/B _12704_/S vssd1 vssd1 vccd1 vccd1 _12704_/X sky130_fd_sc_hd__mux2_1
X_19260_ _19261_/CLK _19260_/D vssd1 vssd1 vccd1 vccd1 _19260_/Q sky130_fd_sc_hd__dfxtp_1
X_16472_ _16538_/A0 _19079_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _19079_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13684_ _19545_/Q _13946_/B vssd1 vssd1 vccd1 vccd1 _13684_/X sky130_fd_sc_hd__or2_1
XFILLER_189_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10896_ _11594_/A1 _18327_/Q _17778_/Q _11605_/S vssd1 vssd1 vccd1 vccd1 _10896_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18211_ _19159_/CLK _18211_/D vssd1 vssd1 vccd1 vccd1 _18211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12635_ _10985_/A _10982_/Y _12634_/X vssd1 vssd1 vccd1 vccd1 _12635_/Y sky130_fd_sc_hd__o21ai_1
X_15423_ _19470_/Q _15498_/S _15422_/Y _15476_/A1 vssd1 vssd1 vccd1 vccd1 _15423_/X
+ sky130_fd_sc_hd__o211a_1
X_19191_ _19625_/CLK _19191_/D vssd1 vssd1 vccd1 vccd1 _19191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18142_ _19627_/CLK _18142_/D vssd1 vssd1 vccd1 vccd1 _18142_/Q sky130_fd_sc_hd__dfxtp_1
X_15354_ _15223_/A _15352_/Y _15353_/X _15416_/A vssd1 vssd1 vccd1 vccd1 _15354_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_200_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12566_ _13165_/C _13167_/B vssd1 vssd1 vccd1 vccd1 _12566_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11517_ _11053_/A _11496_/Y _11502_/Y _11509_/Y _11516_/X vssd1 vssd1 vccd1 vccd1
+ _11517_/X sky130_fd_sc_hd__o32a_4
XFILLER_145_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14305_ _16292_/A0 _18164_/Q _14305_/S vssd1 vssd1 vccd1 vccd1 _18164_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18073_ _19092_/CLK _18073_/D vssd1 vssd1 vccd1 vccd1 _18073_/Q sky130_fd_sc_hd__dfxtp_1
X_15285_ _15304_/A1 _13203_/Y _15285_/A3 _15284_/X vssd1 vssd1 vccd1 vccd1 _15285_/X
+ sky130_fd_sc_hd__a31o_1
X_12497_ _12578_/A _12545_/A vssd1 vssd1 vccd1 vccd1 _12497_/Y sky130_fd_sc_hd__nor2_4
XFILLER_172_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14236_ _18116_/Q _14266_/B vssd1 vssd1 vccd1 vccd1 _14236_/X sky130_fd_sc_hd__or2_1
X_17024_ _17181_/B _17046_/A2 _17023_/X _17376_/A vssd1 vssd1 vccd1 vccd1 _19348_/D
+ sky130_fd_sc_hd__o211a_1
X_11448_ _11219_/A _10235_/B _10834_/B _09039_/B vssd1 vssd1 vccd1 vccd1 _11448_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_144_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14167_ _16892_/A _14167_/B vssd1 vssd1 vccd1 vccd1 _18081_/D sky130_fd_sc_hd__and2_1
XFILLER_113_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11379_ _18639_/Q _18061_/Q _11379_/S vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13118_ _13988_/B vssd1 vssd1 vccd1 vccd1 _13118_/Y sky130_fd_sc_hd__inv_2
X_18975_ _19592_/CLK _18975_/D vssd1 vssd1 vccd1 vccd1 _18975_/Q sky130_fd_sc_hd__dfxtp_1
X_14098_ _17681_/A0 _18038_/Q _14098_/S vssd1 vssd1 vccd1 vccd1 _18038_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13049_ _13863_/B2 _13043_/Y _13048_/X _12712_/S _13045_/X vssd1 vssd1 vccd1 vccd1
+ _13049_/X sky130_fd_sc_hd__o221a_4
X_17926_ _17930_/CLK _17926_/D vssd1 vssd1 vccd1 vccd1 _17926_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1260 _09367_/B vssd1 vssd1 vccd1 vccd1 _09948_/B sky130_fd_sc_hd__buf_8
XFILLER_267_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1271 _14527_/Y vssd1 vssd1 vccd1 vccd1 _14591_/A2 sky130_fd_sc_hd__buf_4
Xfanout1282 _15918_/A2 vssd1 vssd1 vccd1 vccd1 _15906_/A2 sky130_fd_sc_hd__buf_4
X_17857_ _18691_/CLK _17857_/D vssd1 vssd1 vccd1 vccd1 _17857_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_254_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1293 _14591_/B1 vssd1 vssd1 vccd1 vccd1 _14575_/B1 sky130_fd_sc_hd__buf_4
XFILLER_254_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16808_ _16808_/A _16808_/B _16810_/B vssd1 vssd1 vccd1 vccd1 _19291_/D sky130_fd_sc_hd__nor3_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17788_ _19615_/CLK _17788_/D vssd1 vssd1 vccd1 vccd1 _17788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19527_ _19533_/CLK _19527_/D vssd1 vssd1 vccd1 vccd1 _19527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16739_ _19266_/Q _19265_/Q _16739_/C vssd1 vssd1 vccd1 vccd1 _16742_/B sky130_fd_sc_hd__and3_1
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19458_ _19458_/CLK _19458_/D vssd1 vssd1 vccd1 vccd1 _19458_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09211_ _18542_/Q _18417_/Q _10353_/S vssd1 vssd1 vccd1 vccd1 _09211_/X sky130_fd_sc_hd__mux2_1
XFILLER_223_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18409_ _19620_/CLK _18409_/D vssd1 vssd1 vccd1 vccd1 _18409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19389_ _19553_/CLK _19389_/D vssd1 vssd1 vccd1 vccd1 _19389_/Q sky130_fd_sc_hd__dfxtp_1
X_09142_ _11490_/B _09144_/C vssd1 vssd1 vccd1 vccd1 _12598_/B sky130_fd_sc_hd__and2_1
XFILLER_277_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09073_ _15549_/A _17914_/Q _17913_/Q _09073_/D vssd1 vssd1 vccd1 vccd1 _12443_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_148_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09975_ _10275_/S _09973_/X _09974_/X _08967_/S vssd1 vssd1 vccd1 vccd1 _09975_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08926_ _12051_/A _17802_/Q _08932_/A vssd1 vssd1 vccd1 vccd1 _08996_/B sky130_fd_sc_hd__o21bai_2
XFILLER_58_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08857_ _09992_/A vssd1 vssd1 vccd1 vccd1 _08857_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _13647_/A vssd1 vssd1 vccd1 vccd1 _10750_/Y sky130_fd_sc_hd__inv_2
XFILLER_213_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ _09407_/X _09408_/X _09429_/S vssd1 vssd1 vccd1 vccd1 _09409_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10681_ _11143_/A1 _10679_/Y _10680_/X vssd1 vssd1 vccd1 vccd1 _10681_/X sky130_fd_sc_hd__o21a_1
XFILLER_205_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12420_ _12420_/A1 _12432_/A2 _08988_/X _12420_/B1 _18400_/Q vssd1 vssd1 vccd1 vccd1
+ _12421_/B sky130_fd_sc_hd__o32ai_4
XFILLER_185_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12351_ _11695_/B _09991_/A _09649_/X _12432_/B1 _18377_/Q vssd1 vssd1 vccd1 vccd1
+ _12352_/B sky130_fd_sc_hd__o32ai_4
Xclkbuf_leaf_67_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19604_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11302_ _18640_/Q _18062_/Q _11302_/S vssd1 vssd1 vccd1 vccd1 _11302_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15070_ _18554_/Q _16548_/A0 _15070_/S vssd1 vssd1 vccd1 vccd1 _18554_/D sky130_fd_sc_hd__mux2_1
X_12282_ _18089_/Q _12305_/A2 _12305_/B1 _18512_/Q vssd1 vssd1 vccd1 vccd1 _12478_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14021_ _14033_/A1 _13691_/X _14020_/X _14417_/A vssd1 vssd1 vccd1 vccd1 _17975_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_181_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11233_ _18031_/Q _17999_/Q _11247_/S vssd1 vssd1 vccd1 vccd1 _11233_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11164_ _19211_/Q _11482_/A2 _11163_/X _11406_/B2 vssd1 vssd1 vccd1 vccd1 _11164_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_96_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10115_ _10169_/S _10115_/B vssd1 vssd1 vccd1 vccd1 _10115_/X sky130_fd_sc_hd__or2_1
XFILLER_67_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18760_ _18775_/CLK _18760_/D vssd1 vssd1 vccd1 vccd1 _18760_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15972_ _18701_/Q _15953_/B _15976_/B1 _18750_/Q _15976_/C1 vssd1 vssd1 vccd1 vccd1
+ _15972_/X sky130_fd_sc_hd__a221o_1
X_11095_ _11305_/A1 _18150_/Q _18796_/Q _11094_/S vssd1 vssd1 vccd1 vccd1 _11095_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17711_ _17711_/A0 _19637_/Q _17718_/S vssd1 vssd1 vccd1 vccd1 _19637_/D sky130_fd_sc_hd__mux2_1
XFILLER_276_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14923_ _14921_/X _14922_/X _14714_/B vssd1 vssd1 vccd1 vccd1 _14923_/X sky130_fd_sc_hd__a21o_1
X_10046_ _18532_/Q _18407_/Q _10726_/S vssd1 vssd1 vccd1 vccd1 _10046_/X sky130_fd_sc_hd__mux2_1
X_18691_ _18691_/CLK _18691_/D vssd1 vssd1 vccd1 vccd1 _18691_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17642_ _17708_/A0 _19570_/Q _17648_/S vssd1 vssd1 vccd1 vccd1 _19570_/D sky130_fd_sc_hd__mux2_1
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14854_ _19229_/Q _15014_/B _14934_/C _14854_/D vssd1 vssd1 vccd1 vccd1 _14854_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_236_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13805_ _15133_/A _13801_/Y _13804_/X _13869_/B2 vssd1 vssd1 vccd1 vccd1 _13806_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17573_ _17573_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17573_/X sky130_fd_sc_hd__or2_1
XFILLER_205_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11997_ _17764_/Q _17665_/A0 _12019_/S vssd1 vssd1 vccd1 vccd1 _17764_/D sky130_fd_sc_hd__mux2_1
X_14785_ _14785_/A vssd1 vssd1 vccd1 vccd1 _14785_/Y sky130_fd_sc_hd__inv_2
XFILLER_251_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19312_ _19363_/CLK _19312_/D vssd1 vssd1 vccd1 vccd1 _19312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16524_ _16557_/A0 _19130_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _19130_/D sky130_fd_sc_hd__mux2_1
X_13736_ _18125_/Q _13736_/B vssd1 vssd1 vccd1 vccd1 _13737_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10948_ _11332_/B1 _10946_/X _10947_/X vssd1 vssd1 vccd1 vccd1 _11850_/A sky130_fd_sc_hd__o21ai_1
XFILLER_90_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19243_ _19280_/CLK _19243_/D vssd1 vssd1 vccd1 vccd1 _19243_/Q sky130_fd_sc_hd__dfxtp_2
X_16455_ _19063_/Q _16455_/A1 _16457_/S vssd1 vssd1 vccd1 vccd1 _19063_/D sky130_fd_sc_hd__mux2_1
X_13667_ _10754_/A _13912_/A2 _13912_/B1 vssd1 vssd1 vccd1 vccd1 _13667_/Y sky130_fd_sc_hd__a21oi_1
X_10879_ _10877_/X _10878_/X _11127_/S vssd1 vssd1 vccd1 vccd1 _10879_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _18115_/Q _15786_/A2 _15405_/X _15429_/A2 vssd1 vssd1 vccd1 vccd1 _15408_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_19174_ _19206_/CLK _19174_/D vssd1 vssd1 vccd1 vccd1 _19174_/Q sky130_fd_sc_hd__dfxtp_1
X_12618_ _13148_/B _13148_/C _13148_/A vssd1 vssd1 vccd1 vccd1 _13188_/B sky130_fd_sc_hd__a21oi_2
X_16386_ _16486_/A0 _18997_/Q _16388_/S vssd1 vssd1 vccd1 vccd1 _18997_/D sky130_fd_sc_hd__mux2_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _13861_/A _14147_/C _13892_/B1 vssd1 vssd1 vccd1 vccd1 _13598_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18125_ _19448_/CLK _18125_/D vssd1 vssd1 vccd1 vccd1 _18125_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_247_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12549_ _17823_/Q _13105_/B _12547_/X _12540_/X _12548_/X vssd1 vssd1 vccd1 vccd1
+ _12549_/X sky130_fd_sc_hd__o221a_1
X_15337_ _15335_/X _15364_/A vssd1 vssd1 vccd1 vccd1 _15365_/D sky130_fd_sc_hd__and2b_1
XFILLER_129_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18056_ _19636_/CLK _18056_/D vssd1 vssd1 vccd1 vccd1 _18056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _18197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15268_ _15365_/A _15268_/B vssd1 vssd1 vccd1 vccd1 _15268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_133_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17007_ _19340_/Q _17009_/B vssd1 vssd1 vccd1 vccd1 _17007_/X sky130_fd_sc_hd__or2_1
XFILLER_160_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14219_ _18281_/Q _14267_/A2 _14218_/X _16052_/A vssd1 vssd1 vccd1 vccd1 _18107_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15199_ _15199_/A _15199_/B vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__xnor2_1
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout508 _17499_/A2 vssd1 vssd1 vccd1 vccd1 _17517_/B sky130_fd_sc_hd__clkbuf_2
Xfanout519 _17244_/B vssd1 vssd1 vccd1 vccd1 _17241_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_58_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09760_ _11084_/S _09755_/X _09759_/X vssd1 vssd1 vccd1 vccd1 _09768_/A sky130_fd_sc_hd__o21ai_1
XFILLER_113_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18958_ _19118_/CLK _18958_/D vssd1 vssd1 vccd1 vccd1 _18958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17909_ _17982_/CLK _17909_/D vssd1 vssd1 vccd1 vccd1 _17909_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09691_ _09690_/A _09673_/Y _09690_/Y _09350_/S vssd1 vssd1 vccd1 vccd1 _09691_/X
+ sky130_fd_sc_hd__a211o_1
X_18889_ _19216_/CLK _18889_/D vssd1 vssd1 vccd1 vccd1 _18889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_273_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1090 _17662_/A0 vssd1 vssd1 vccd1 vccd1 _16595_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09125_ _11465_/A1 _19629_/Q _18918_/Q _11455_/S vssd1 vssd1 vccd1 vccd1 _09125_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09056_ _11055_/B2 _08985_/X _09105_/A _11518_/B2 vssd1 vssd1 vccd1 vccd1 _15332_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09958_ _09708_/A _09953_/X _09957_/X _09958_/C1 vssd1 vssd1 vccd1 vccd1 _09958_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_185_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18973_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_277_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _17793_/Q _17792_/Q vssd1 vssd1 vccd1 vccd1 _08929_/B sky130_fd_sc_hd__or2_4
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_114_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19285_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _11189_/A _09887_/X _09888_/X _11198_/S vssd1 vssd1 vccd1 vccd1 _09889_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11920_ _11926_/A1 _11939_/A1 _11803_/B _11935_/B1 input215/X vssd1 vssd1 vccd1 vccd1
+ _11920_/X sky130_fd_sc_hd__a32o_4
XFILLER_46_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_402 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_413 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11851_ _11859_/B _11816_/X _11791_/Y _11801_/A vssd1 vssd1 vccd1 vccd1 _11851_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_424 _11774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_435 _12550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10802_ _19120_/Q _19152_/Q _11605_/S vssd1 vssd1 vccd1 vccd1 _10802_/X sky130_fd_sc_hd__mux2_1
XANTENNA_446 _14008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_457 _18576_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _14576_/A _14570_/B vssd1 vssd1 vccd1 vccd1 _18393_/D sky130_fd_sc_hd__or2_1
XANTENNA_468 _18397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11782_ _11816_/A _11782_/B vssd1 vssd1 vccd1 vccd1 _11803_/B sky130_fd_sc_hd__nor2_8
XANTENNA_479 input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13521_ _19508_/Q _13781_/A2 _13947_/B1 _13520_/X vssd1 vssd1 vccd1 vccd1 _13521_/X
+ sky130_fd_sc_hd__o211a_1
X_10733_ _18616_/Q _18187_/Q _10744_/S vssd1 vssd1 vccd1 vccd1 _10733_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16240_ _11452_/B _18855_/Q _16255_/S vssd1 vssd1 vccd1 vccd1 _18855_/D sky130_fd_sc_hd__mux2_1
X_13452_ _19506_/Q _13781_/A2 _13947_/B1 _13451_/X vssd1 vssd1 vccd1 vccd1 _13452_/X
+ sky130_fd_sc_hd__o211a_1
X_10664_ _10660_/X _10663_/X _11601_/A vssd1 vssd1 vccd1 vccd1 _10664_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12403_ _12430_/A _12403_/B vssd1 vssd1 vccd1 vccd1 _12403_/Y sky130_fd_sc_hd__nand2_1
XFILLER_167_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16171_ _17701_/A0 _18788_/Q _16192_/S vssd1 vssd1 vccd1 vccd1 _18788_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13383_ _13758_/A _13369_/Y _13956_/B1 vssd1 vssd1 vccd1 vccd1 _13383_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10595_ _10589_/S _10590_/Y _10594_/Y _11602_/C1 vssd1 vssd1 vccd1 vccd1 _10595_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12334_ _08929_/X _12333_/X _12325_/X vssd1 vssd1 vccd1 vccd1 _12334_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15122_ _15118_/A _15118_/B _17124_/A _15123_/B vssd1 vssd1 vccd1 vccd1 _15122_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15053_ _18537_/Q _17664_/A0 _15076_/S vssd1 vssd1 vccd1 vccd1 _18537_/D sky130_fd_sc_hd__mux2_1
X_12265_ _12837_/A _12265_/B vssd1 vssd1 vccd1 vccd1 _12265_/Y sky130_fd_sc_hd__nand2_4
XFILLER_154_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14004_ _14004_/A _14004_/B vssd1 vssd1 vccd1 vccd1 _14004_/Y sky130_fd_sc_hd__nand2_1
X_11216_ _17967_/Q _11216_/A2 _11216_/B1 vssd1 vssd1 vccd1 vccd1 _11216_/X sky130_fd_sc_hd__a21o_1
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12196_ _17862_/Q _12194_/B _12195_/Y vssd1 vssd1 vccd1 vccd1 _17862_/D sky130_fd_sc_hd__o21a_1
X_18812_ _19619_/CLK _18812_/D vssd1 vssd1 vccd1 vccd1 _18812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11147_ _18642_/Q _18064_/Q _11147_/S vssd1 vssd1 vccd1 vccd1 _11147_/X sky130_fd_sc_hd__mux2_1
XFILLER_268_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18743_ _18746_/CLK _18743_/D vssd1 vssd1 vccd1 vccd1 _18743_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15955_ _15953_/A _15955_/B vssd1 vssd1 vccd1 vccd1 _15955_/Y sky130_fd_sc_hd__nand2b_1
X_11078_ _11559_/S1 _11077_/X _11076_/X _11084_/S vssd1 vssd1 vccd1 vccd1 _11078_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput160 dout1[58] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_hd__buf_2
XFILLER_236_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput171 irq[0] vssd1 vssd1 vccd1 vccd1 input171/X sky130_fd_sc_hd__clkbuf_4
XFILLER_264_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14906_ input56/X input91/X _14947_/S vssd1 vssd1 vccd1 vccd1 _14907_/A sky130_fd_sc_hd__mux2_2
Xinput182 irq[5] vssd1 vssd1 vccd1 vccd1 _15086_/C sky130_fd_sc_hd__buf_2
X_10029_ _19035_/Q _19003_/Q _11609_/S vssd1 vssd1 vccd1 vccd1 _10029_/X sky130_fd_sc_hd__mux2_1
X_18674_ _18715_/CLK _18674_/D vssd1 vssd1 vccd1 vccd1 _18674_/Q sky130_fd_sc_hd__dfxtp_1
Xinput193 localMemory_wb_adr_i[12] vssd1 vssd1 vccd1 vccd1 input193/X sky130_fd_sc_hd__clkbuf_2
XFILLER_270_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15886_ _18671_/Q _15949_/A2 _15885_/X _15904_/C1 vssd1 vssd1 vccd1 vccd1 _18671_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _17625_/A _17658_/A vssd1 vssd1 vccd1 vccd1 _17625_/Y sky130_fd_sc_hd__nand2_8
XFILLER_52_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14837_ _14833_/Y _14836_/X _14950_/B1 vssd1 vssd1 vccd1 vccd1 _14837_/Y sky130_fd_sc_hd__a21oi_4
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17556_ _17556_/A _17589_/B vssd1 vssd1 vccd1 vccd1 _17556_/X sky130_fd_sc_hd__and2_4
XFILLER_189_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14768_ _17798_/Q _14911_/B vssd1 vssd1 vccd1 vccd1 _14768_/X sky130_fd_sc_hd__or2_1
XFILLER_17_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16507_ _16507_/A0 _19113_/Q _16524_/S vssd1 vssd1 vccd1 vccd1 _19113_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13719_ _19448_/Q _13949_/A2 _13717_/X _13718_/X _13949_/C1 vssd1 vssd1 vccd1 vccd1
+ _13719_/X sky130_fd_sc_hd__o221a_2
XFILLER_177_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17487_ _18120_/Q _17539_/C1 _17485_/X _17486_/X vssd1 vssd1 vccd1 vccd1 _17487_/X
+ sky130_fd_sc_hd__a22o_1
X_14699_ _14875_/B1 _14695_/X _14698_/Y _14928_/B1 vssd1 vssd1 vccd1 vccd1 _14700_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_220_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19226_ _19226_/CLK _19226_/D vssd1 vssd1 vccd1 vccd1 _19226_/Q sky130_fd_sc_hd__dfxtp_1
X_16438_ _19046_/Q _09105_/A _16457_/S vssd1 vssd1 vccd1 vccd1 _19046_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19157_ _19157_/CLK _19157_/D vssd1 vssd1 vccd1 vccd1 _19157_/Q sky130_fd_sc_hd__dfxtp_1
X_16369_ _16535_/A0 _18980_/Q _16390_/S vssd1 vssd1 vccd1 vccd1 _18980_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18108_ _18778_/CLK _18108_/D vssd1 vssd1 vccd1 vccd1 _18108_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_258_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19088_ _19226_/CLK _19088_/D vssd1 vssd1 vccd1 vccd1 _19088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18039_ _19154_/CLK _18039_/D vssd1 vssd1 vccd1 vccd1 _18039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_278_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09812_ _11279_/B1 _09811_/X _09796_/Y _09791_/X vssd1 vssd1 vccd1 vccd1 _09812_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09743_ _09859_/A _09743_/B vssd1 vssd1 vccd1 vccd1 _11790_/C sky130_fd_sc_hd__nor2_1
XFILLER_28_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09674_ _18536_/Q _18411_/Q _18020_/Q _17988_/Q _09688_/S _10266_/S1 vssd1 vssd1
+ vccd1 vccd1 _09674_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09108_ _10623_/A _09108_/B _09853_/S _09108_/D vssd1 vssd1 vccd1 vccd1 _09108_/X
+ sky130_fd_sc_hd__or4_4
X_10380_ _11550_/A vssd1 vssd1 vccd1 vccd1 _10380_/Y sky130_fd_sc_hd__inv_2
X_09039_ _11556_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _09042_/A sky130_fd_sc_hd__or2_2
XFILLER_191_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12050_ _17900_/Q _12052_/A2 _12049_/X _13257_/A vssd1 vssd1 vccd1 vccd1 _17802_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11001_ _11469_/A1 _19572_/Q _11386_/S _19604_/Q _11001_/C1 vssd1 vssd1 vccd1 vccd1
+ _11001_/X sky130_fd_sc_hd__o221a_1
Xfanout1804 _15039_/A vssd1 vssd1 vccd1 vccd1 _14427_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1815 _17380_/A vssd1 vssd1 vccd1 vccd1 _17354_/A sky130_fd_sc_hd__buf_4
Xfanout1826 _17336_/A vssd1 vssd1 vccd1 vccd1 _17350_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_120_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1837 _13987_/C1 vssd1 vssd1 vccd1 vccd1 _14417_/A sky130_fd_sc_hd__buf_4
Xfanout1848 _17342_/A vssd1 vssd1 vccd1 vccd1 _17346_/A sky130_fd_sc_hd__buf_4
Xfanout850 _10792_/A2 vssd1 vssd1 vccd1 vccd1 _17713_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_266_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout861 _10609_/X vssd1 vssd1 vccd1 vccd1 _16615_/A0 sky130_fd_sc_hd__buf_4
XFILLER_265_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1859 fanout1863/X vssd1 vssd1 vccd1 vccd1 _14205_/A sky130_fd_sc_hd__buf_4
XFILLER_277_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout872 _10238_/X vssd1 vssd1 vccd1 vccd1 _10239_/B sky130_fd_sc_hd__buf_4
XFILLER_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout883 _12813_/S vssd1 vssd1 vccd1 vccd1 _12818_/S sky130_fd_sc_hd__buf_4
Xfanout894 _12936_/S vssd1 vssd1 vccd1 vccd1 _13039_/S sky130_fd_sc_hd__buf_2
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ _15782_/A1 _15739_/X _15782_/B1 vssd1 vssd1 vccd1 vccd1 _15740_/X sky130_fd_sc_hd__a21o_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _12952_/A vssd1 vssd1 vccd1 vccd1 _12952_/Y sky130_fd_sc_hd__inv_2
XFILLER_252_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11903_ _11903_/A _11903_/B vssd1 vssd1 vccd1 vccd1 _11904_/B sky130_fd_sc_hd__nor2_8
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _15671_/A _15671_/B vssd1 vssd1 vccd1 vccd1 _15672_/B sky130_fd_sc_hd__nor2_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _18566_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12883_ _12883_/A vssd1 vssd1 vccd1 vccd1 _12883_/Y sky130_fd_sc_hd__inv_2
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_221 _18640_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 _18390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _11737_/X _15118_/A _15117_/A _17794_/Q _15116_/B vssd1 vssd1 vccd1 vccd1
+ _17410_/X sky130_fd_sc_hd__a221o_1
XANTENNA_243 _18380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _16548_/A0 _18429_/Q _14622_/S vssd1 vssd1 vccd1 vccd1 _18429_/D sky130_fd_sc_hd__mux2_1
XANTENNA_254 _15087_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11834_ _14141_/B _11834_/B vssd1 vssd1 vccd1 vccd1 _11834_/Y sky130_fd_sc_hd__nand2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _19399_/CLK _18390_/D vssd1 vssd1 vccd1 vccd1 _18390_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 input225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 input240/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _19468_/Q _17583_/A _17377_/S vssd1 vssd1 vccd1 vccd1 _17342_/B sky130_fd_sc_hd__mux2_1
XANTENNA_287 _11899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_298 _18735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11765_ _18583_/Q _14349_/B _11770_/B1 _13622_/B vssd1 vssd1 vccd1 vccd1 _11765_/X
+ sky130_fd_sc_hd__a22o_4
X_14553_ _18385_/Q _14559_/A2 _14559_/B1 input13/X vssd1 vssd1 vccd1 vccd1 _14554_/B
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_82_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19206_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _13682_/B2 _13493_/X _13494_/Y _13503_/Y vssd1 vssd1 vccd1 vccd1 _14008_/B
+ sky130_fd_sc_hd__o2bb2a_4
X_10716_ _12320_/A _11135_/S _11181_/B1 _10715_/Y vssd1 vssd1 vccd1 vccd1 _10753_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_158_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17272_ _18118_/Q _17219_/A _17478_/A _17310_/B vssd1 vssd1 vccd1 vccd1 _17272_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14484_ _18336_/Q _17688_/A0 _14485_/S vssd1 vssd1 vccd1 vccd1 _18336_/D sky130_fd_sc_hd__mux2_1
X_11696_ _11687_/Y _11692_/X _11694_/Y _11695_/X _12461_/A vssd1 vssd1 vccd1 vccd1
+ _11696_/X sky130_fd_sc_hd__o2111a_1
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19640_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19011_ _19213_/CLK _19011_/D vssd1 vssd1 vccd1 vccd1 _19011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16223_ _16455_/A1 _18839_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _18839_/D sky130_fd_sc_hd__mux2_1
X_13435_ _13747_/B2 _13423_/X _13424_/Y _13434_/Y vssd1 vssd1 vccd1 vccd1 _14004_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ _18071_/Q _10816_/A2 _10646_/X _10643_/S vssd1 vssd1 vccd1 vccd1 _10647_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_228_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16154_ _16154_/A _16154_/B _16154_/C vssd1 vssd1 vccd1 vccd1 _18776_/D sky130_fd_sc_hd__and3_1
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13366_ _13937_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _13366_/X sky130_fd_sc_hd__or2_1
X_10578_ _11112_/A _10570_/X _10569_/X _10653_/C1 vssd1 vssd1 vccd1 vccd1 _10578_/X
+ sky130_fd_sc_hd__a211o_1
X_15105_ _14158_/A _14158_/B _14158_/C _15328_/B vssd1 vssd1 vccd1 vccd1 _15124_/C
+ sky130_fd_sc_hd__o31ai_4
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12317_ _12442_/C _13260_/B vssd1 vssd1 vccd1 vccd1 _12317_/X sky130_fd_sc_hd__or2_1
X_13297_ _19244_/Q _13495_/A2 _13495_/B1 _19276_/Q vssd1 vssd1 vccd1 vccd1 _13297_/X
+ sky130_fd_sc_hd__a22o_1
X_16085_ _18745_/Q _16093_/B vssd1 vssd1 vccd1 vccd1 _16085_/Y sky130_fd_sc_hd__nand2_1
XFILLER_269_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15036_ _18525_/Q _12269_/A _15037_/S vssd1 vssd1 vccd1 vccd1 _18525_/D sky130_fd_sc_hd__mux2_1
X_12248_ _17881_/Q _17882_/Q _12248_/C vssd1 vssd1 vccd1 vccd1 _12253_/C sky130_fd_sc_hd__and3_2
XFILLER_268_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12179_ _12187_/A _12184_/C vssd1 vssd1 vccd1 vccd1 _12179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_284_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16987_ _19330_/Q _17043_/B vssd1 vssd1 vccd1 vccd1 _16987_/X sky130_fd_sc_hd__or2_1
XFILLER_256_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18726_ _18734_/CLK _18726_/D vssd1 vssd1 vccd1 vccd1 _18726_/Q sky130_fd_sc_hd__dfxtp_1
X_15938_ input5/X input280/X _15947_/S vssd1 vssd1 vccd1 vccd1 _15938_/X sky130_fd_sc_hd__mux2_1
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18657_ _19586_/CLK _18657_/D vssd1 vssd1 vccd1 vccd1 _18657_/Q sky130_fd_sc_hd__dfxtp_4
X_15869_ _15869_/A _15905_/B _15908_/C vssd1 vssd1 vccd1 vccd1 _15869_/X sky130_fd_sc_hd__and3_1
XFILLER_236_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17608_ _19545_/Q _17624_/A2 _17607_/X _17368_/A vssd1 vssd1 vccd1 vccd1 _19545_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09390_ _19107_/Q _19139_/Q _10353_/S vssd1 vssd1 vccd1 vccd1 _09390_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18588_ _19450_/CLK _18588_/D vssd1 vssd1 vccd1 vccd1 _18588_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17539_ _18591_/Q _17538_/A _17538_/Y _17539_/C1 vssd1 vssd1 vccd1 vccd1 _17539_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_225_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19209_ _19216_/CLK _19209_/D vssd1 vssd1 vccd1 vccd1 _19209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput420 _18490_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[19] sky130_fd_sc_hd__buf_4
XFILLER_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput431 _18500_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[29] sky130_fd_sc_hd__buf_4
Xoutput442 _18529_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_stall_o sky130_fd_sc_hd__buf_4
XFILLER_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput453 _18113_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[12] sky130_fd_sc_hd__buf_4
Xoutput464 _18123_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[22] sky130_fd_sc_hd__buf_4
Xoutput475 _18104_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[3] sky130_fd_sc_hd__buf_4
XFILLER_160_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput486 _11957_/X vssd1 vssd1 vccd1 vccd1 wmask0[2] sky130_fd_sc_hd__buf_4
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09726_ _09976_/A1 _09724_/X _09725_/X _08967_/S vssd1 vssd1 vccd1 vccd1 _09726_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_216_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09657_ input119/X input154/X _09657_/S vssd1 vssd1 vccd1 vccd1 _09657_/X sky130_fd_sc_hd__mux2_8
XFILLER_83_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09588_ _18444_/Q _18345_/Q _10362_/S vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__mux2_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11550_ _11550_/A _11550_/B vssd1 vssd1 vccd1 vccd1 _13812_/A sky130_fd_sc_hd__nor2_8
XFILLER_184_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ _08901_/A _18229_/Q _10500_/S _18964_/Q _10033_/S vssd1 vssd1 vccd1 vccd1
+ _10501_/X sky130_fd_sc_hd__o221a_1
XFILLER_184_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11481_ _11481_/A _18791_/Q _11481_/C vssd1 vssd1 vccd1 vccd1 _11481_/X sky130_fd_sc_hd__and3_1
XFILLER_168_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13220_ _13289_/A _13218_/Y _13219_/X _11751_/A _13916_/A vssd1 vssd1 vccd1 vccd1
+ _13220_/X sky130_fd_sc_hd__o32a_1
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10432_ _19061_/Q _19029_/Q _10656_/S vssd1 vssd1 vccd1 vccd1 _10432_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13151_ _12685_/X _12737_/X _13354_/A vssd1 vssd1 vccd1 vccd1 _13152_/A sky130_fd_sc_hd__mux2_1
X_10363_ _10361_/X _10362_/X _10371_/S vssd1 vssd1 vccd1 vccd1 _10363_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ _17827_/Q _12098_/B _12101_/Y vssd1 vssd1 vccd1 vccd1 _17827_/D sky130_fd_sc_hd__o21a_1
XFILLER_152_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13082_ _13083_/B _13083_/C _13083_/A vssd1 vssd1 vccd1 vccd1 _13126_/B sky130_fd_sc_hd__a21o_1
X_10294_ _10294_/A1 _18161_/Q _18807_/Q _10299_/S vssd1 vssd1 vccd1 vccd1 _10294_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16910_ _16848_/S _17936_/Q _16909_/X vssd1 vssd1 vccd1 vccd1 _17169_/B sky130_fd_sc_hd__o21a_4
X_12033_ _17794_/Q _12051_/B vssd1 vssd1 vccd1 vccd1 _12033_/X sky130_fd_sc_hd__or2_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1601 _08887_/Y vssd1 vssd1 vccd1 vccd1 _11663_/A sky130_fd_sc_hd__clkbuf_16
Xfanout1612 _16137_/B vssd1 vssd1 vccd1 vccd1 _16139_/B sky130_fd_sc_hd__buf_4
X_17890_ _17901_/CLK _17890_/D vssd1 vssd1 vccd1 vccd1 _17890_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1623 _12432_/A2 vssd1 vssd1 vccd1 vccd1 _09232_/A sky130_fd_sc_hd__buf_6
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1634 _08864_/X vssd1 vssd1 vccd1 vccd1 _15082_/A sky130_fd_sc_hd__buf_6
X_16841_ _17048_/A _17217_/A vssd1 vssd1 vccd1 vccd1 _17316_/A sky130_fd_sc_hd__or2_4
Xfanout1645 _10817_/A1 vssd1 vssd1 vccd1 vccd1 _10662_/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1656 _09873_/A1 vssd1 vssd1 vccd1 vccd1 _10219_/A1 sky130_fd_sc_hd__buf_8
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1667 _08849_/Y vssd1 vssd1 vccd1 vccd1 _10030_/C1 sky130_fd_sc_hd__clkbuf_16
XFILLER_120_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout680 _13247_/A2 vssd1 vssd1 vccd1 vccd1 _13951_/A2 sky130_fd_sc_hd__buf_8
Xfanout1678 _11584_/A1 vssd1 vssd1 vccd1 vccd1 _11305_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_92_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1689 _12468_/B vssd1 vssd1 vccd1 vccd1 _10262_/A1 sky130_fd_sc_hd__buf_6
X_19560_ _19592_/CLK _19560_/D vssd1 vssd1 vccd1 vccd1 _19560_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout691 _13655_/C1 vssd1 vssd1 vccd1 vccd1 _13949_/C1 sky130_fd_sc_hd__buf_4
XFILLER_120_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16772_ _19278_/Q _16775_/C _16780_/B1 vssd1 vssd1 vccd1 vccd1 _16772_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_247_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13984_ _17957_/Q _14004_/A vssd1 vssd1 vccd1 vccd1 _13984_/X sky130_fd_sc_hd__or2_1
XFILLER_19_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18511_ _19321_/CLK _18511_/D vssd1 vssd1 vccd1 vccd1 _18511_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15723_ _15723_/A _15723_/B vssd1 vssd1 vccd1 vccd1 _15724_/A sky130_fd_sc_hd__nor2_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _12813_/X _12818_/X _12935_/S vssd1 vssd1 vccd1 vccd1 _12935_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19491_ _19525_/CLK _19491_/D vssd1 vssd1 vccd1 vccd1 _19491_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18442_ _19621_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _19480_/Q _15653_/Y _15716_/S vssd1 vssd1 vccd1 vccd1 _15654_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _13757_/A _13978_/B _12847_/X vssd1 vssd1 vccd1 vccd1 _12866_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_261_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _17664_/A0 _18412_/Q _14628_/S vssd1 vssd1 vccd1 vccd1 _18412_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11817_ _11865_/A _11816_/X _11815_/Y vssd1 vssd1 vccd1 vccd1 _11818_/C sky130_fd_sc_hd__a21oi_4
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _19399_/CLK _18373_/D vssd1 vssd1 vccd1 vccd1 _18373_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15585_ _15789_/B1 _15583_/Y _15584_/Y _12322_/Y vssd1 vssd1 vccd1 vccd1 _15585_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12797_ _12696_/X _12687_/X _12818_/S vssd1 vssd1 vccd1 vccd1 _12797_/X sky130_fd_sc_hd__mux2_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17324_ _17565_/B _17377_/S _17323_/Y _17330_/A vssd1 vssd1 vccd1 vccd1 _19459_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _14596_/A _14536_/B vssd1 vssd1 vccd1 vccd1 _18376_/D sky130_fd_sc_hd__or2_1
X_11748_ _13148_/A _11748_/B vssd1 vssd1 vccd1 vccd1 _13147_/A sky130_fd_sc_hd__xnor2_4
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ _17255_/A _17255_/B vssd1 vssd1 vccd1 vccd1 _19435_/D sky130_fd_sc_hd__nor2_1
X_14467_ _18319_/Q _17671_/A0 _14483_/S vssd1 vssd1 vccd1 vccd1 _18319_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ _12626_/B _11679_/B vssd1 vssd1 vccd1 vccd1 _13402_/B sky130_fd_sc_hd__xnor2_4
X_16206_ _17703_/A0 _18822_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _18822_/D sky130_fd_sc_hd__mux2_1
X_13418_ _13411_/A _14155_/B _13417_/Y _11293_/B vssd1 vssd1 vccd1 vccd1 _13418_/X
+ sky130_fd_sc_hd__o22a_1
X_17186_ _17285_/A _17186_/B vssd1 vssd1 vccd1 vccd1 _19413_/D sky130_fd_sc_hd__nor2_1
X_14398_ _17705_/A0 _18249_/Q _14415_/S vssd1 vssd1 vccd1 vccd1 _18249_/D sky130_fd_sc_hd__mux2_1
X_16137_ _18771_/Q _16137_/B vssd1 vssd1 vccd1 vccd1 _16137_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13349_ _13366_/B _13349_/B vssd1 vssd1 vccd1 vccd1 _13349_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16068_ _11981_/B _16069_/A _16054_/A _18741_/Q vssd1 vssd1 vccd1 vccd1 _16068_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15019_ _18508_/Q input208/X _16627_/S vssd1 vssd1 vccd1 vccd1 _18508_/D sky130_fd_sc_hd__mux2_1
X_08890_ _17894_/Q _17893_/Q _09070_/D _12439_/A vssd1 vssd1 vccd1 vccd1 _08890_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_229_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09511_ _11190_/A1 _19560_/Q _09724_/S _19592_/Q _09723_/S vssd1 vssd1 vccd1 vccd1
+ _09511_/X sky130_fd_sc_hd__o221a_1
X_18709_ _18761_/CLK _18709_/D vssd1 vssd1 vccd1 vccd1 _18709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09442_ _10263_/A1 _18211_/Q _09671_/S _18946_/Q _10266_/S1 vssd1 vssd1 vccd1 vccd1
+ _09442_/X sky130_fd_sc_hd__o221a_1
XFILLER_25_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _18602_/Q _18173_/Q _09966_/S vssd1 vssd1 vccd1 vccd1 _09373_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput294 _11910_/X vssd1 vssd1 vccd1 vccd1 addr1[0] sky130_fd_sc_hd__buf_4
XFILLER_248_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09709_ _09708_/A _09706_/X _09708_/Y _09958_/C1 vssd1 vssd1 vccd1 vccd1 _09709_/X
+ sky130_fd_sc_hd__o211a_1
X_10981_ _18120_/Q _10980_/Y _11135_/S vssd1 vssd1 vccd1 vccd1 _10985_/B sky130_fd_sc_hd__mux2_2
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12720_ _11061_/B _11445_/B _12721_/S vssd1 vssd1 vccd1 vccd1 _12720_/X sky130_fd_sc_hd__mux2_4
XFILLER_74_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12651_ _13763_/A _12650_/X _12649_/X vssd1 vssd1 vccd1 vccd1 _12651_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11602_ _11601_/A _11599_/X _11601_/Y _11602_/C1 vssd1 vssd1 vccd1 vccd1 _11602_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_169_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12582_ _12582_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _12582_/X sky130_fd_sc_hd__or2_4
X_15370_ _19436_/Q _15124_/B _15354_/X _15369_/X _17166_/A vssd1 vssd1 vccd1 vccd1
+ _15370_/X sky130_fd_sc_hd__o221a_1
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14321_ _18178_/Q _17705_/A0 _14338_/S vssd1 vssd1 vccd1 vccd1 _18178_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11533_ _13533_/A _11675_/B _11673_/A _11060_/Y vssd1 vssd1 vccd1 vccd1 _11534_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_183_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17040_ _17205_/B _17046_/A2 _17039_/X _17374_/A vssd1 vssd1 vccd1 vccd1 _19356_/D
+ sky130_fd_sc_hd__o211a_1
X_11464_ _11465_/A1 _19566_/Q _11462_/S _19598_/Q _11464_/C1 vssd1 vssd1 vccd1 vccd1
+ _11464_/X sky130_fd_sc_hd__o221a_1
XFILLER_183_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14252_ _14252_/A _14252_/B vssd1 vssd1 vccd1 vccd1 _14252_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10415_ _11411_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10415_/Y sky130_fd_sc_hd__nor2_1
X_13203_ _13203_/A vssd1 vssd1 vccd1 vccd1 _13203_/Y sky130_fd_sc_hd__inv_2
X_11395_ _11481_/A _19176_/Q _11395_/C vssd1 vssd1 vccd1 vccd1 _11395_/X sky130_fd_sc_hd__and3_1
X_14183_ _16153_/D _14183_/B vssd1 vssd1 vccd1 vccd1 _18089_/D sky130_fd_sc_hd__and2_1
XFILLER_174_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10346_ _10344_/X _10345_/X _10346_/S vssd1 vssd1 vccd1 vccd1 _10346_/X sky130_fd_sc_hd__mux2_1
X_13134_ _12930_/X _12935_/X _13134_/S vssd1 vssd1 vccd1 vccd1 _13414_/B sky130_fd_sc_hd__mux2_1
X_18991_ _19611_/CLK _18991_/D vssd1 vssd1 vccd1 vccd1 _18991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17942_ _19231_/CLK _17942_/D vssd1 vssd1 vccd1 vccd1 _17942_/Q sky130_fd_sc_hd__dfxtp_1
X_13065_ _19528_/Q _13277_/S _13243_/B1 vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__o21a_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10277_ _18044_/Q _18012_/Q _10299_/S vssd1 vssd1 vccd1 vccd1 _10277_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1420 _11384_/B vssd1 vssd1 vccd1 vccd1 _11386_/S sky130_fd_sc_hd__buf_4
XFILLER_266_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12016_ _17783_/Q _16551_/A0 _12022_/S vssd1 vssd1 vccd1 vccd1 _17783_/D sky130_fd_sc_hd__mux2_1
Xfanout1431 _10009_/A vssd1 vssd1 vccd1 vccd1 _10326_/A sky130_fd_sc_hd__buf_12
X_17873_ _19324_/CLK _17873_/D vssd1 vssd1 vccd1 vccd1 _17873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1442 _11002_/C1 vssd1 vssd1 vccd1 vccd1 _09935_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_238_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1453 _10337_/S1 vssd1 vssd1 vccd1 vccd1 _10266_/S1 sky130_fd_sc_hd__buf_6
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1464 fanout1469/X vssd1 vssd1 vccd1 vccd1 _11360_/B2 sky130_fd_sc_hd__buf_6
X_19612_ _19612_/CLK _19612_/D vssd1 vssd1 vccd1 vccd1 _19612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_266_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16824_ _16824_/A _16981_/B vssd1 vssd1 vccd1 vccd1 _17048_/A sky130_fd_sc_hd__nand2_1
Xfanout1475 fanout1525/X vssd1 vssd1 vccd1 vccd1 _10511_/S sky130_fd_sc_hd__buf_6
XFILLER_281_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1486 _10496_/B vssd1 vssd1 vccd1 vccd1 _10500_/S sky130_fd_sc_hd__buf_6
XFILLER_226_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1497 _10290_/S vssd1 vssd1 vccd1 vccd1 _09704_/S sky130_fd_sc_hd__buf_6
XFILLER_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19543_ _19543_/CLK _19543_/D vssd1 vssd1 vccd1 vccd1 _19543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16755_ _16768_/A _16755_/B _16759_/C vssd1 vssd1 vccd1 vccd1 _19271_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13967_ _13259_/X _13958_/X _13961_/X _13966_/X vssd1 vssd1 vccd1 vccd1 _13967_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_62_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15706_ _15746_/C _15706_/B vssd1 vssd1 vccd1 vccd1 _15706_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12918_ _12917_/X _15866_/A _12918_/S vssd1 vssd1 vccd1 vccd1 _12918_/X sky130_fd_sc_hd__mux2_1
XFILLER_235_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19474_ _19540_/CLK _19474_/D vssd1 vssd1 vccd1 vccd1 _19474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16686_ _16740_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16686_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13898_ _12444_/X _13897_/Y _13889_/X _13322_/Y vssd1 vssd1 vccd1 vccd1 _13899_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18425_ _19636_/CLK _18425_/D vssd1 vssd1 vccd1 vccd1 _18425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_261_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15637_ _15744_/A _15687_/A vssd1 vssd1 vccd1 vccd1 _15686_/A sky130_fd_sc_hd__xnor2_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _19458_/Q _12768_/A _13165_/C _13925_/S vssd1 vssd1 vccd1 vccd1 _12849_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_222_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18356_ _19634_/CLK _18356_/D vssd1 vssd1 vccd1 vccd1 _18356_/Q sky130_fd_sc_hd__dfxtp_1
X_15568_ _15568_/A _15568_/B vssd1 vssd1 vccd1 vccd1 _15570_/A sky130_fd_sc_hd__nand2_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17307_ _19453_/Q _17307_/B vssd1 vssd1 vccd1 vccd1 _17307_/Y sky130_fd_sc_hd__nand2_1
X_14519_ _17721_/A0 _18369_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _18369_/D sky130_fd_sc_hd__mux2_1
XFILLER_202_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18287_ _19448_/CLK _18287_/D vssd1 vssd1 vccd1 vccd1 _18287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15499_ _17219_/A _15498_/X _15499_/B1 vssd1 vssd1 vccd1 vccd1 _15499_/X sky130_fd_sc_hd__a21o_1
X_17238_ _19430_/Q _17256_/B vssd1 vssd1 vccd1 vccd1 _17238_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17169_ _17214_/A _17169_/B vssd1 vssd1 vccd1 vccd1 _17473_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ _09991_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__nor2_1
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ _17794_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08942_/Y sky130_fd_sc_hd__nor2_2
XFILLER_103_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08873_ _10513_/S _09494_/A _12755_/A _17900_/Q vssd1 vssd1 vccd1 vccd1 _08875_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ _18243_/Q _18818_/Q _18446_/Q _18347_/Q _09428_/B2 _09978_/A1 vssd1 vssd1
+ vccd1 vccd1 _09426_/B sky130_fd_sc_hd__mux4_1
XFILLER_252_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _11001_/C1 _09355_/X _09354_/X _11478_/S vssd1 vssd1 vccd1 vccd1 _09360_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_139_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19490_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09287_ _18603_/Q _18174_/Q _09302_/S vssd1 vssd1 vccd1 vccd1 _09287_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10200_ _10198_/X _10199_/X _10200_/S vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ _11488_/A _11837_/A vssd1 vssd1 vccd1 vccd1 _11180_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10131_ _10225_/S _10130_/X _10129_/X _11046_/S1 vssd1 vssd1 vccd1 vccd1 _10131_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_279_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10062_ _18101_/Q _10061_/X _11441_/B vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__mux2_8
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14870_ _18488_/Q _15001_/A2 _14869_/Y _16803_/A vssd1 vssd1 vccd1 vccd1 _18488_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13821_ _17850_/Q _13821_/B vssd1 vssd1 vccd1 vccd1 _13821_/Y sky130_fd_sc_hd__nor2_1
XFILLER_235_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16540_ _16540_/A0 _19145_/Q _16557_/S vssd1 vssd1 vccd1 vccd1 _19145_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13752_ _19353_/Q _13883_/A2 _13883_/B1 _19481_/Q _13883_/C1 vssd1 vssd1 vccd1 vccd1
+ _13752_/X sky130_fd_sc_hd__a221o_1
XFILLER_232_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10964_ _11360_/A1 _19214_/Q _19182_/Q _11340_/B2 vssd1 vssd1 vccd1 vccd1 _10964_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12703_ _12601_/B _12658_/B _12704_/S vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__mux2_1
X_16471_ _16471_/A0 _19078_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _19078_/D sky130_fd_sc_hd__mux2_1
XFILLER_231_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ _19319_/Q _13174_/A _13722_/B1 _13682_/X vssd1 vssd1 vccd1 vccd1 _13683_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10895_ _11594_/A1 _19606_/Q _19574_/Q _11605_/S vssd1 vssd1 vccd1 vccd1 _10895_/X
+ sky130_fd_sc_hd__a22o_1
X_18210_ _18445_/CLK _18210_/D vssd1 vssd1 vccd1 vccd1 _18210_/Q sky130_fd_sc_hd__dfxtp_1
X_15422_ _15498_/S _15422_/B vssd1 vssd1 vccd1 vccd1 _15422_/Y sky130_fd_sc_hd__nand2_1
XPHY_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19190_ _19623_/CLK _19190_/D vssd1 vssd1 vccd1 vccd1 _19190_/Q sky130_fd_sc_hd__dfxtp_1
X_12634_ _13568_/A _12634_/B vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__or2_1
XFILLER_70_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18141_ _19626_/CLK _18141_/D vssd1 vssd1 vccd1 vccd1 _18141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15353_ _18574_/Q _15388_/C vssd1 vssd1 vccd1 vccd1 _15353_/X sky130_fd_sc_hd__or2_1
X_12565_ _12584_/A _13167_/B vssd1 vssd1 vccd1 vccd1 _12565_/X sky130_fd_sc_hd__or2_1
XFILLER_129_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14304_ _16622_/A0 _18163_/Q _14304_/S vssd1 vssd1 vccd1 vccd1 _18163_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11516_ _11511_/Y _11515_/Y _11516_/B1 vssd1 vssd1 vccd1 vccd1 _11516_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18072_ _19611_/CLK _18072_/D vssd1 vssd1 vccd1 vccd1 _18072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15284_ _15284_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _15284_/X sky130_fd_sc_hd__and2_1
X_12496_ _12548_/A _12554_/B vssd1 vssd1 vccd1 vccd1 _12545_/A sky130_fd_sc_hd__nand2b_4
XFILLER_8_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17023_ _19348_/Q _17041_/B vssd1 vssd1 vccd1 vccd1 _17023_/X sky130_fd_sc_hd__or2_1
XFILLER_144_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14235_ _18289_/Q _14261_/A2 _14234_/X _14451_/B vssd1 vssd1 vccd1 vccd1 _18115_/D
+ sky130_fd_sc_hd__o211a_1
X_11447_ _17964_/Q _11447_/A2 _09899_/X vssd1 vssd1 vccd1 vccd1 _11447_/X sky130_fd_sc_hd__a21o_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11378_ _19080_/Q _11462_/S _11377_/X _11464_/C1 vssd1 vssd1 vccd1 vccd1 _11378_/X
+ sky130_fd_sc_hd__o211a_1
X_14166_ _18694_/Q _18081_/Q _14200_/S vssd1 vssd1 vccd1 vccd1 _14167_/B sky130_fd_sc_hd__mux2_1
XFILLER_171_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10329_ _10334_/A1 _17785_/Q _09181_/S _18334_/Q vssd1 vssd1 vccd1 vccd1 _10329_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_252_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13117_ _13115_/B2 _13102_/X _13105_/Y _13116_/Y vssd1 vssd1 vccd1 vccd1 _13988_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_180_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14097_ _17680_/A0 _18037_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _18037_/D sky130_fd_sc_hd__mux2_1
X_18974_ _19114_/CLK _18974_/D vssd1 vssd1 vccd1 vccd1 _18974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13048_ _13390_/S _13047_/Y _13197_/B1 vssd1 vssd1 vccd1 vccd1 _13048_/X sky130_fd_sc_hd__a21o_1
X_17925_ _17930_/CLK _17925_/D vssd1 vssd1 vccd1 vccd1 _17925_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1250 _08930_/Y vssd1 vssd1 vccd1 vccd1 _11447_/A2 sky130_fd_sc_hd__buf_4
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1261 _13237_/B1 vssd1 vssd1 vccd1 vccd1 _09367_/B sky130_fd_sc_hd__buf_6
X_17856_ _19306_/CLK _17856_/D vssd1 vssd1 vccd1 vccd1 _17856_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1272 _12277_/B vssd1 vssd1 vccd1 vccd1 _12305_/A2 sky130_fd_sc_hd__buf_8
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1283 _15918_/A2 vssd1 vssd1 vccd1 vccd1 _15948_/A2 sky130_fd_sc_hd__buf_4
XFILLER_254_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1294 _14528_/X vssd1 vssd1 vccd1 vccd1 _14591_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_226_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16807_ _19291_/Q _19290_/Q _16807_/C vssd1 vssd1 vccd1 vccd1 _16810_/B sky130_fd_sc_hd__and3_2
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17787_ _19615_/CLK _17787_/D vssd1 vssd1 vccd1 vccd1 _17787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14999_ _15009_/A1 _18272_/Q _14998_/Y _11712_/A vssd1 vssd1 vccd1 vccd1 _14999_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16738_ _19265_/Q _16739_/C _16737_/Y vssd1 vssd1 vccd1 vccd1 _19265_/D sky130_fd_sc_hd__o21a_1
XFILLER_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19526_ _19526_/CLK _19526_/D vssd1 vssd1 vccd1 vccd1 _19526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19457_ _19522_/CLK _19457_/D vssd1 vssd1 vccd1 vccd1 _19457_/Q sky130_fd_sc_hd__dfxtp_2
X_16669_ _19244_/Q _16670_/C _16668_/Y vssd1 vssd1 vccd1 vccd1 _19244_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09210_ _18317_/Q _17768_/Q _10353_/S vssd1 vssd1 vccd1 vccd1 _09210_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18408_ _19047_/CLK _18408_/D vssd1 vssd1 vccd1 vccd1 _18408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19388_ _19553_/CLK _19388_/D vssd1 vssd1 vccd1 vccd1 _19388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09141_ _09141_/A _11103_/A vssd1 vssd1 vccd1 vccd1 _11592_/S sky130_fd_sc_hd__nor2_1
X_18339_ _19625_/CLK _18339_/D vssd1 vssd1 vccd1 vccd1 _18339_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_277_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09072_ _17901_/Q _12264_/B vssd1 vssd1 vccd1 vccd1 _12740_/B sky130_fd_sc_hd__or2_4
XFILLER_129_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _11497_/A1 _18205_/Q _09952_/S _18940_/Q _09972_/S vssd1 vssd1 vccd1 vccd1
+ _09974_/X sky130_fd_sc_hd__o221a_1
XFILLER_130_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08925_ _12051_/A _17802_/Q _08932_/A vssd1 vssd1 vccd1 vccd1 _08995_/B sky130_fd_sc_hd__o21ba_4
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08856_ _17792_/Q vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__inv_2
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09408_ _10294_/A1 _18314_/Q _17765_/Q _09428_/B2 vssd1 vssd1 vccd1 vccd1 _09408_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10680_ _17974_/Q _16820_/A3 _11216_/B1 vssd1 vssd1 vccd1 vccd1 _10680_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09339_ _11404_/A1 _17766_/Q _09344_/S _18315_/Q _10250_/S vssd1 vssd1 vccd1 vccd1
+ _09339_/X sky130_fd_sc_hd__o221a_1
XFILLER_187_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ _17891_/Q _12382_/A _12349_/Y _12350_/C1 vssd1 vssd1 vccd1 vccd1 _17891_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_275_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11301_ _19081_/Q _11302_/S _11300_/X _11311_/C1 vssd1 vssd1 vccd1 vccd1 _11301_/X
+ sky130_fd_sc_hd__o211a_1
X_12281_ _18094_/Q _12305_/A2 _12305_/B1 _18517_/Q vssd1 vssd1 vccd1 vccd1 _12285_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14020_ _17975_/Q _14020_/B vssd1 vssd1 vccd1 vccd1 _14020_/X sky130_fd_sc_hd__or2_1
XFILLER_153_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11232_ _18422_/Q _11224_/B _11231_/X _11567_/S vssd1 vssd1 vccd1 vccd1 _11232_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11163_ _11173_/S _19179_/Q _11171_/S vssd1 vssd1 vccd1 vccd1 _11163_/X sky130_fd_sc_hd__and3_1
XFILLER_121_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19626_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10114_ _10112_/X _10113_/X _10335_/S vssd1 vssd1 vccd1 vccd1 _10115_/B sky130_fd_sc_hd__mux2_1
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15971_ _18701_/Q _15977_/A2 _15970_/X _14181_/A vssd1 vssd1 vccd1 vccd1 _18701_/D
+ sky130_fd_sc_hd__o211a_1
X_11094_ _18860_/Q _18892_/Q _11094_/S vssd1 vssd1 vccd1 vccd1 _11094_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17710_ _17710_/A0 _19636_/Q _17719_/S vssd1 vssd1 vccd1 vccd1 _19636_/D sky130_fd_sc_hd__mux2_1
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10045_ _18307_/Q _17758_/Q _11617_/S vssd1 vssd1 vccd1 vccd1 _10045_/X sky130_fd_sc_hd__mux2_1
X_14922_ _15003_/A1 _13691_/X _15003_/B1 _18649_/Q _15003_/C1 vssd1 vssd1 vccd1 vccd1
+ _14922_/X sky130_fd_sc_hd__a221o_1
X_18690_ _18691_/CLK _18690_/D vssd1 vssd1 vccd1 vccd1 _18690_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _17641_/A0 _19569_/Q _17657_/S vssd1 vssd1 vccd1 vccd1 _19569_/D sky130_fd_sc_hd__mux2_1
XFILLER_263_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14853_ _14238_/A _14893_/S _14851_/X _14852_/X vssd1 vssd1 vccd1 vccd1 _14853_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_264_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _13837_/B _13804_/B vssd1 vssd1 vccd1 vccd1 _13804_/X sky130_fd_sc_hd__or2_2
XFILLER_263_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17572_ _19528_/Q _17561_/B _17588_/B1 _17571_/X vssd1 vssd1 vccd1 vccd1 _19528_/D
+ sky130_fd_sc_hd__o211a_1
X_14784_ input106/X input78/X _14784_/S vssd1 vssd1 vccd1 vccd1 _14785_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11996_ _17763_/Q _17664_/A0 _12019_/S vssd1 vssd1 vccd1 vccd1 _17763_/D sky130_fd_sc_hd__mux2_1
X_19311_ _19324_/CLK _19311_/D vssd1 vssd1 vccd1 vccd1 _19311_/Q sky130_fd_sc_hd__dfxtp_1
X_16523_ _16622_/A0 _19129_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _19129_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13735_ _18125_/Q _13736_/B vssd1 vssd1 vccd1 vccd1 _13802_/C sky130_fd_sc_hd__and2_1
X_10947_ _10532_/A _16545_/A0 _11800_/B vssd1 vssd1 vccd1 vccd1 _10947_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19242_ _19276_/CLK _19242_/D vssd1 vssd1 vccd1 vccd1 _19242_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_220_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16454_ _19062_/Q _16619_/A0 _16454_/S vssd1 vssd1 vccd1 vccd1 _19062_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13666_ _13761_/B _14149_/B vssd1 vssd1 vccd1 vccd1 _13666_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ _11596_/A1 _18614_/Q _18185_/Q _10815_/B vssd1 vssd1 vccd1 vccd1 _10878_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15405_ _15404_/B _13399_/X _15133_/B _15404_/Y vssd1 vssd1 vccd1 vccd1 _15405_/X
+ sky130_fd_sc_hd__a31o_1
X_19173_ _19594_/CLK _19173_/D vssd1 vssd1 vccd1 vccd1 _19173_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _13127_/A _13126_/A _12616_/X _12615_/A _12612_/Y vssd1 vssd1 vccd1 vccd1
+ _13148_/C sky130_fd_sc_hd__o221a_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _17684_/A0 _18996_/Q _16385_/S vssd1 vssd1 vccd1 vccd1 _18996_/D sky130_fd_sc_hd__mux2_1
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _13597_/A _13597_/B vssd1 vssd1 vccd1 vccd1 _14147_/C sky130_fd_sc_hd__xnor2_1
X_18124_ _19444_/CLK _18124_/D vssd1 vssd1 vccd1 vccd1 _18124_/Q sky130_fd_sc_hd__dfxtp_4
X_15336_ _15335_/B _15336_/B vssd1 vssd1 vccd1 vccd1 _15364_/A sky130_fd_sc_hd__nand2b_2
XFILLER_184_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12548_ _12548_/A _12768_/B vssd1 vssd1 vccd1 vccd1 _12548_/X sky130_fd_sc_hd__or2_4
XFILLER_247_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18055_ _19138_/CLK _18055_/D vssd1 vssd1 vccd1 vccd1 _18055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15267_ _15365_/A _15268_/B vssd1 vssd1 vccd1 vccd1 _15267_/X sky130_fd_sc_hd__or2_1
X_12479_ _16821_/A _08841_/Y _12478_/Y vssd1 vssd1 vccd1 vccd1 _12502_/A sky130_fd_sc_hd__a21oi_1
XANTENNA_2 _18197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17006_ _17581_/A _17044_/A2 _17005_/X _17346_/A vssd1 vssd1 vccd1 vccd1 _19339_/D
+ sky130_fd_sc_hd__o211a_1
X_14218_ _18107_/Q _14244_/B vssd1 vssd1 vccd1 vccd1 _14218_/X sky130_fd_sc_hd__or2_1
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15198_ _15199_/A _15199_/B vssd1 vssd1 vccd1 vccd1 _15198_/X sky130_fd_sc_hd__or2_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14149_ _14149_/A _14149_/B _14149_/C _14149_/D vssd1 vssd1 vccd1 vccd1 _14151_/C
+ sky130_fd_sc_hd__or4_2
Xfanout509 _17499_/A2 vssd1 vssd1 vccd1 vccd1 _17547_/B sky130_fd_sc_hd__buf_6
XFILLER_141_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18957_ _19604_/CLK _18957_/D vssd1 vssd1 vccd1 vccd1 _18957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17908_ _17982_/CLK _17908_/D vssd1 vssd1 vccd1 vccd1 _17908_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09690_ _09690_/A _09690_/B vssd1 vssd1 vccd1 vccd1 _09690_/Y sky130_fd_sc_hd__nor2_1
XFILLER_273_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18888_ _19208_/CLK _18888_/D vssd1 vssd1 vccd1 vccd1 _18888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1080 _09980_/A2 vssd1 vssd1 vccd1 vccd1 _17693_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_254_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1091 _16529_/A0 vssd1 vssd1 vccd1 vccd1 _17662_/A0 sky130_fd_sc_hd__buf_2
X_17839_ _19310_/CLK _17839_/D vssd1 vssd1 vccd1 vccd1 _17839_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19509_ _19521_/CLK _19509_/D vssd1 vssd1 vccd1 vccd1 _19509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09124_ _12466_/A0 _09120_/X _09123_/X _11459_/B1 vssd1 vssd1 vccd1 vccd1 _09124_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09055_ _08958_/A _09055_/B _09055_/C vssd1 vssd1 vccd1 vccd1 _09055_/X sky130_fd_sc_hd__and3b_1
XFILLER_190_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09957_ _09954_/X _09955_/X _09956_/X _10742_/A1 _10301_/S vssd1 vssd1 vccd1 vccd1
+ _09957_/X sky130_fd_sc_hd__a221o_1
XFILLER_89_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ _08816_/A _17791_/Q _17790_/Q vssd1 vssd1 vccd1 vccd1 _08940_/B sky130_fd_sc_hd__nand3b_4
XFILLER_246_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09888_ _08901_/A _18206_/Q _10054_/S _18941_/Q _10033_/S vssd1 vssd1 vccd1 vccd1
+ _09888_/X sky130_fd_sc_hd__o221a_1
XFILLER_218_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08839_ _12442_/A vssd1 vssd1 vccd1 vccd1 _15307_/A sky130_fd_sc_hd__inv_2
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_403 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _11850_/A _11864_/B vssd1 vssd1 vccd1 vccd1 _11850_/X sky130_fd_sc_hd__or2_4
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_414 _10609_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_425 _11822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_154_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19433_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_436 _13978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_447 _13527_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801_ _18069_/Q _10816_/A2 _10800_/X _11611_/S vssd1 vssd1 vccd1 vccd1 _10801_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_458 _18567_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11781_ _15039_/B _11780_/X _11726_/B vssd1 vssd1 vccd1 vccd1 _11781_/X sky130_fd_sc_hd__a21o_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_469 _18401_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13520_ _19540_/Q _13946_/B vssd1 vssd1 vccd1 vccd1 _13520_/X sky130_fd_sc_hd__or2_1
XFILLER_242_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10732_ _18258_/Q _18833_/Q _10744_/S vssd1 vssd1 vccd1 vccd1 _10732_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13451_ _19538_/Q _13946_/B vssd1 vssd1 vccd1 vccd1 _13451_/X sky130_fd_sc_hd__or2_1
X_10663_ _10661_/X _10662_/X _10663_/S vssd1 vssd1 vccd1 vccd1 _10663_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12402_ _12420_/A1 _09236_/A _09571_/X _12429_/B1 _18394_/Q vssd1 vssd1 vccd1 vccd1
+ _12403_/B sky130_fd_sc_hd__o32ai_2
XFILLER_185_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16170_ _16203_/A0 _18787_/Q _16189_/S vssd1 vssd1 vccd1 vccd1 _18787_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10594_ _11601_/A _10594_/B vssd1 vssd1 vccd1 vccd1 _10594_/Y sky130_fd_sc_hd__nor2_1
X_13382_ _13637_/A _14002_/B _13369_/Y vssd1 vssd1 vccd1 vccd1 _13382_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15121_ _08882_/B _15117_/A _15120_/Y _17461_/A2 _17559_/B vssd1 vssd1 vccd1 vccd1
+ _17124_/A sky130_fd_sc_hd__o311a_4
X_12333_ _15047_/B _12333_/B _12333_/C _12333_/D vssd1 vssd1 vccd1 vccd1 _12333_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_127_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15052_ _18536_/Q _17696_/A0 _15076_/S vssd1 vssd1 vccd1 vccd1 _18536_/D sky130_fd_sc_hd__mux2_1
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12264_ _12264_/A _12264_/B _12837_/A vssd1 vssd1 vccd1 vccd1 _12264_/X sky130_fd_sc_hd__and3_2
XFILLER_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14003_ _17966_/Q _14028_/A _14002_/Y _14181_/A vssd1 vssd1 vccd1 vccd1 _17966_/D
+ sky130_fd_sc_hd__o211a_1
X_11215_ _13468_/S _11215_/B vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__nor2_4
X_12195_ _16752_/A _12200_/C vssd1 vssd1 vccd1 vccd1 _12195_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18811_ _18875_/CLK _18811_/D vssd1 vssd1 vccd1 vccd1 _18811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_268_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _19083_/Q _11147_/S _11145_/X _11156_/C1 vssd1 vssd1 vccd1 vccd1 _11146_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18742_ _18749_/CLK _18742_/D vssd1 vssd1 vccd1 vccd1 _18742_/Q sky130_fd_sc_hd__dfxtp_2
X_15954_ _18731_/Q _15954_/B _15955_/B vssd1 vssd1 vccd1 vccd1 _15954_/X sky130_fd_sc_hd__and3_1
X_11077_ _18033_/Q _18001_/Q _11094_/S vssd1 vssd1 vccd1 vccd1 _11077_/X sky130_fd_sc_hd__mux2_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput150 dout1[49] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_hd__clkbuf_2
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput161 dout1[59] vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_hd__buf_2
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905_ _15006_/A1 _14904_/X _15006_/B1 vssd1 vssd1 vccd1 vccd1 _14905_/Y sky130_fd_sc_hd__o21ai_2
Xinput172 irq[10] vssd1 vssd1 vccd1 vccd1 _15091_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10028_ _10026_/X _10027_/Y _09141_/A vssd1 vssd1 vccd1 vccd1 _10028_/X sky130_fd_sc_hd__a21o_1
X_18673_ _18683_/CLK _18673_/D vssd1 vssd1 vccd1 vccd1 _18673_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15885_ _18670_/Q _15906_/A2 _15948_/C1 _15884_/X vssd1 vssd1 vccd1 vccd1 _15885_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput183 irq[6] vssd1 vssd1 vccd1 vccd1 input183/X sky130_fd_sc_hd__buf_2
Xinput194 localMemory_wb_adr_i[13] vssd1 vssd1 vccd1 vccd1 input194/X sky130_fd_sc_hd__clkbuf_2
XFILLER_236_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ _15009_/A1 _18270_/Q _14835_/Y _14918_/B1 vssd1 vssd1 vccd1 vccd1 _14836_/X
+ sky130_fd_sc_hd__a31o_2
X_17624_ _19553_/Q _17624_/A2 _17591_/X _17214_/B _17623_/X vssd1 vssd1 vccd1 vccd1
+ _19553_/D sky130_fd_sc_hd__o221a_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _17555_/A _17555_/B _17591_/C vssd1 vssd1 vccd1 vccd1 _17555_/X sky130_fd_sc_hd__or3_1
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14767_ _18478_/Q _14720_/A _14766_/Y _12243_/A vssd1 vssd1 vccd1 vccd1 _18478_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11979_ _18737_/Q _18734_/Q _11979_/C vssd1 vssd1 vccd1 vccd1 _15954_/B sky130_fd_sc_hd__nor3_4
XFILLER_204_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16506_ _16539_/A0 _19112_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _19112_/D sky130_fd_sc_hd__mux2_1
XFILLER_205_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13718_ _19416_/Q _13948_/A2 _13948_/B1 vssd1 vssd1 vccd1 vccd1 _13718_/X sky130_fd_sc_hd__a21o_1
XFILLER_205_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17486_ _18581_/Q _17544_/A _08883_/A vssd1 vssd1 vccd1 vccd1 _17486_/X sky130_fd_sc_hd__o21a_1
X_14698_ _14718_/A _14698_/B vssd1 vssd1 vccd1 vccd1 _14698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19225_ _19225_/CLK _19225_/D vssd1 vssd1 vccd1 vccd1 _19225_/Q sky130_fd_sc_hd__dfxtp_1
X_16437_ _19045_/Q _16602_/A0 _16457_/S vssd1 vssd1 vccd1 vccd1 _19045_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ _17845_/Q _13846_/B _12548_/X vssd1 vssd1 vccd1 vccd1 _13649_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19156_ _19620_/CLK _19156_/D vssd1 vssd1 vccd1 vccd1 _19156_/Q sky130_fd_sc_hd__dfxtp_1
X_16368_ _16501_/A0 _18979_/Q _16390_/S vssd1 vssd1 vccd1 vccd1 _18979_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18107_ _18741_/CLK _18107_/D vssd1 vssd1 vccd1 vccd1 _18107_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15319_ _19466_/Q _19400_/Q vssd1 vssd1 vccd1 vccd1 _15319_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19087_ _19618_/CLK _19087_/D vssd1 vssd1 vccd1 vccd1 _19087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16299_ _17697_/A0 _18912_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _18912_/D sky130_fd_sc_hd__mux2_1
XFILLER_274_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18038_ _19645_/CLK _18038_/D vssd1 vssd1 vccd1 vccd1 _18038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09811_ _11622_/C1 _09805_/X _09808_/X _09810_/X vssd1 vssd1 vccd1 vccd1 _09811_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_259_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09742_ _17955_/Q _11216_/A2 _08947_/X _17923_/Q _09741_/X vssd1 vssd1 vccd1 vccd1
+ _09743_/B sky130_fd_sc_hd__a221o_4
XFILLER_228_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09673_ _11173_/S _09671_/X _09672_/X vssd1 vssd1 vccd1 vccd1 _09673_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09107_ _09108_/D _10633_/A _10838_/B _09107_/D vssd1 vssd1 vccd1 vccd1 _11790_/B
+ sky130_fd_sc_hd__and4b_4
XFILLER_109_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09038_ _10309_/A _11219_/A _09037_/X _09019_/Y vssd1 vssd1 vccd1 vccd1 _09038_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11000_ _11001_/C1 _10999_/X _10998_/X _11478_/S vssd1 vssd1 vccd1 vccd1 _11000_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_104_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1805 fanout1870/X vssd1 vssd1 vccd1 vccd1 _15039_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_77_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1816 _17366_/A vssd1 vssd1 vccd1 vccd1 _17368_/A sky130_fd_sc_hd__buf_4
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1827 _17336_/A vssd1 vssd1 vccd1 vccd1 _17469_/C1 sky130_fd_sc_hd__buf_4
XFILLER_278_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout840 _10989_/X vssd1 vssd1 vccd1 vccd1 _17710_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout1838 _14179_/A vssd1 vssd1 vccd1 vccd1 _14037_/C1 sky130_fd_sc_hd__buf_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1849 _13987_/C1 vssd1 vssd1 vccd1 vccd1 _17342_/A sky130_fd_sc_hd__buf_4
Xfanout851 _10792_/A2 vssd1 vssd1 vccd1 vccd1 _16580_/A0 sky130_fd_sc_hd__clkbuf_2
Xfanout862 _10609_/X vssd1 vssd1 vccd1 vccd1 _17682_/A0 sky130_fd_sc_hd__buf_4
Xfanout873 _10166_/X vssd1 vssd1 vccd1 vccd1 _16621_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_284_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout884 _12796_/S vssd1 vssd1 vccd1 vccd1 _12813_/S sky130_fd_sc_hd__buf_4
XFILLER_265_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout895 _12602_/A vssd1 vssd1 vccd1 vccd1 _12936_/S sky130_fd_sc_hd__clkbuf_4
X_12951_ _13314_/S _12990_/B _12745_/X vssd1 vssd1 vccd1 vccd1 _12952_/A sky130_fd_sc_hd__a21boi_1
XFILLER_86_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _11828_/X _11875_/A _11875_/Y _11829_/Y _11901_/X vssd1 vssd1 vccd1 vccd1
+ _11903_/B sky130_fd_sc_hd__o221a_4
X_15670_ _19481_/Q _19415_/Q vssd1 vssd1 vccd1 vccd1 _15671_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 _14036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12882_ _12830_/X _12881_/X _13134_/S vssd1 vssd1 vccd1 vccd1 _12883_/A sky130_fd_sc_hd__mux2_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 _18568_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _18655_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _17680_/A0 _18428_/Q _14631_/S vssd1 vssd1 vccd1 vccd1 _18428_/D sky130_fd_sc_hd__mux2_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 _18392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11833_ _11833_/A vssd1 vssd1 vccd1 vccd1 _11833_/Y sky130_fd_sc_hd__clkinv_2
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_244 _18382_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _15087_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_266 input226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17559_/A _17340_/B vssd1 vssd1 vccd1 vccd1 _19467_/D sky130_fd_sc_hd__and2_1
XANTENNA_277 input241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14576_/A _14552_/B vssd1 vssd1 vccd1 vccd1 _18384_/D sky130_fd_sc_hd__or2_1
XFILLER_186_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_288 _11920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _18582_/Q _14349_/B _11769_/B1 _13611_/B vssd1 vssd1 vccd1 vccd1 _11764_/X
+ sky130_fd_sc_hd__a22o_4
XANTENNA_299 _18735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _19313_/Q _13174_/A _13722_/B1 _13496_/X _13502_/X vssd1 vssd1 vccd1 vccd1
+ _13503_/Y sky130_fd_sc_hd__a2111oi_2
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _11103_/A _11864_/A vssd1 vssd1 vccd1 vccd1 _10715_/Y sky130_fd_sc_hd__nor2_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _19441_/Q _17310_/B vssd1 vssd1 vccd1 vccd1 _17271_/Y sky130_fd_sc_hd__nand2_1
X_14483_ _18335_/Q _16488_/A0 _14483_/S vssd1 vssd1 vccd1 vccd1 _18335_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11695_ _18268_/Q _11695_/B vssd1 vssd1 vccd1 vccd1 _11695_/X sky130_fd_sc_hd__or2_2
X_19010_ _19614_/CLK _19010_/D vssd1 vssd1 vccd1 vccd1 _19010_/Q sky130_fd_sc_hd__dfxtp_1
X_16222_ _16619_/A0 _18838_/Q _16222_/S vssd1 vssd1 vccd1 vccd1 _18838_/D sky130_fd_sc_hd__mux2_1
X_13434_ _19311_/Q _13754_/A2 _13426_/X _13427_/X _13433_/X vssd1 vssd1 vccd1 vccd1
+ _13434_/Y sky130_fd_sc_hd__a2111oi_2
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10646_ _18649_/Q _10650_/S vssd1 vssd1 vccd1 vccd1 _10646_/X sky130_fd_sc_hd__or2_1
XFILLER_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ _18776_/Q _18775_/Q _18774_/Q _16153_/D vssd1 vssd1 vccd1 vccd1 _16154_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_158_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13365_ _13937_/A _13365_/B vssd1 vssd1 vccd1 vccd1 _13365_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_wb_clk_i clkbuf_leaf_79_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19203_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_166_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10577_ _11112_/A _10575_/X _10576_/X _10653_/C1 vssd1 vssd1 vccd1 vccd1 _10577_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_177_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ _18778_/Q _18777_/Q vssd1 vssd1 vccd1 vccd1 _15104_/X sky130_fd_sc_hd__or2_2
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12316_ _12442_/C _13260_/B vssd1 vssd1 vccd1 vccd1 _15303_/B sky130_fd_sc_hd__nor2_4
X_16084_ _16096_/A1 _16083_/Y _17725_/C1 vssd1 vssd1 vccd1 vccd1 _18744_/D sky130_fd_sc_hd__a21oi_1
XFILLER_6_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13296_ _17835_/Q _13844_/A2 _13844_/B1 _17867_/Q vssd1 vssd1 vccd1 vccd1 _13296_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15035_ _18524_/Q _12269_/B _15037_/S vssd1 vssd1 vccd1 vccd1 _18524_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12247_ _17881_/Q _12248_/C _17882_/Q vssd1 vssd1 vccd1 vccd1 _12249_/B sky130_fd_sc_hd__a21oi_1
XFILLER_244_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12178_ _17856_/Q _12178_/B vssd1 vssd1 vccd1 vccd1 _12184_/C sky130_fd_sc_hd__and2_2
XFILLER_268_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11129_ _11112_/A _11124_/X _11128_/X vssd1 vssd1 vccd1 vccd1 _11131_/C sky130_fd_sc_hd__a21oi_1
XFILLER_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16986_ _17123_/B _17044_/A2 _16985_/X _17328_/A vssd1 vssd1 vccd1 vccd1 _19329_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_284_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18725_ _18775_/CLK _18725_/D vssd1 vssd1 vccd1 vccd1 _18725_/Q sky130_fd_sc_hd__dfxtp_4
X_15937_ _18688_/Q _15943_/A2 _15936_/X _15946_/C1 vssd1 vssd1 vccd1 vccd1 _18688_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15868_ _18665_/Q _15910_/A2 _15866_/X _15867_/X _15910_/C1 vssd1 vssd1 vccd1 vccd1
+ _18665_/D sky130_fd_sc_hd__o221a_1
X_18656_ _19076_/CLK _18656_/D vssd1 vssd1 vccd1 vccd1 _18656_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_209_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14819_ _12459_/X _14000_/B _14683_/X _18639_/Q vssd1 vssd1 vccd1 vccd1 _14819_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_17607_ _19488_/Q _15085_/X _17556_/A _17190_/B _17556_/X vssd1 vssd1 vccd1 vccd1
+ _17607_/X sky130_fd_sc_hd__a221o_1
XFILLER_92_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15799_ _15797_/Y _15798_/X _15800_/A2 vssd1 vssd1 vccd1 vccd1 _15799_/Y sky130_fd_sc_hd__o21ai_1
X_18587_ _19448_/CLK _18587_/D vssd1 vssd1 vccd1 vccd1 _18587_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_225_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17538_ _17538_/A _17538_/B vssd1 vssd1 vccd1 vccd1 _17538_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17469_ _19505_/Q _17547_/B _17467_/X _17468_/Y _17469_/C1 vssd1 vssd1 vccd1 vccd1
+ _19505_/D sky130_fd_sc_hd__o221a_1
XFILLER_193_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19208_ _19208_/CLK _19208_/D vssd1 vssd1 vccd1 vccd1 _19208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19139_ _19636_/CLK _19139_/D vssd1 vssd1 vccd1 vccd1 _19139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput410 _18471_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[0] sky130_fd_sc_hd__buf_4
Xoutput421 _18472_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[1] sky130_fd_sc_hd__buf_4
XFILLER_218_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput432 _18473_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[2] sky130_fd_sc_hd__buf_4
XFILLER_172_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput443 _08883_/Y vssd1 vssd1 vccd1 vccd1 probe_env[0] sky130_fd_sc_hd__buf_4
XFILLER_271_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput454 _18114_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[13] sky130_fd_sc_hd__buf_4
Xoutput465 _18124_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[23] sky130_fd_sc_hd__buf_4
Xoutput476 _14214_/A vssd1 vssd1 vccd1 vccd1 probe_programCounter[4] sky130_fd_sc_hd__buf_4
XFILLER_232_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput487 _11959_/X vssd1 vssd1 vccd1 vccd1 wmask0[3] sky130_fd_sc_hd__buf_4
XFILLER_102_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09725_ _11190_/A1 _18208_/Q _09724_/S _18943_/Q _09723_/S vssd1 vssd1 vccd1 vccd1
+ _09725_/X sky130_fd_sc_hd__o221a_1
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09656_ _09012_/A _09232_/A _09655_/X _09656_/B1 _18401_/Q vssd1 vssd1 vccd1 vccd1
+ _10234_/B sky130_fd_sc_hd__o32a_1
XFILLER_43_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09587_ _10746_/S _09586_/X _09585_/X _08895_/A vssd1 vssd1 vccd1 vccd1 _09587_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10500_ _19092_/Q _18996_/Q _10500_/S vssd1 vssd1 vccd1 vccd1 _10500_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11480_ _18855_/Q _11481_/C _11479_/X _11480_/C1 vssd1 vssd1 vccd1 vccd1 _11480_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10431_ _08904_/A _10425_/X _10428_/X _10430_/X vssd1 vssd1 vccd1 vccd1 _10431_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13150_ _13224_/B _13149_/X _13147_/Y _12442_/C vssd1 vssd1 vccd1 vccd1 _13150_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_192_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10362_ _18621_/Q _18192_/Q _10362_/S vssd1 vssd1 vccd1 vccd1 _10362_/X sky130_fd_sc_hd__mux2_1
X_12101_ _12107_/A _12106_/C vssd1 vssd1 vccd1 vccd1 _12101_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10293_ _18871_/Q _10290_/S _10293_/B1 vssd1 vssd1 vccd1 vccd1 _10293_/X sky130_fd_sc_hd__o21a_1
X_13081_ _13081_/A _13349_/B vssd1 vssd1 vccd1 vccd1 _13081_/X sky130_fd_sc_hd__and2_1
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12032_ _17891_/Q _12035_/B _12031_/X _12350_/C1 vssd1 vssd1 vccd1 vccd1 _17793_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1602 _08887_/Y vssd1 vssd1 vccd1 vccd1 _11918_/A2 sky130_fd_sc_hd__buf_4
Xfanout1613 _16095_/B vssd1 vssd1 vccd1 vccd1 _16137_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1624 _08987_/Y vssd1 vssd1 vccd1 vccd1 _12432_/A2 sky130_fd_sc_hd__buf_4
Xfanout1635 _12420_/A1 vssd1 vssd1 vccd1 vccd1 _11695_/B sky130_fd_sc_hd__buf_6
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16840_ _16981_/A _16840_/B _16981_/B vssd1 vssd1 vccd1 vccd1 _17555_/A sky130_fd_sc_hd__nand3b_1
Xfanout1646 _09873_/A1 vssd1 vssd1 vccd1 vccd1 _10817_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout1657 _09873_/A1 vssd1 vssd1 vccd1 vccd1 _10354_/A1 sky130_fd_sc_hd__buf_4
XFILLER_120_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1668 _15481_/A vssd1 vssd1 vccd1 vccd1 _11602_/C1 sky130_fd_sc_hd__buf_6
Xfanout670 _11824_/A vssd1 vssd1 vccd1 vccd1 _14141_/B sky130_fd_sc_hd__buf_8
Xfanout681 _12565_/X vssd1 vssd1 vccd1 vccd1 _13247_/A2 sky130_fd_sc_hd__buf_6
Xfanout1679 _10625_/A1 vssd1 vssd1 vccd1 vccd1 _11584_/A1 sky130_fd_sc_hd__buf_8
XFILLER_120_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16771_ _16776_/A _16771_/B _16775_/C vssd1 vssd1 vccd1 vccd1 _19277_/D sky130_fd_sc_hd__nor3_1
XFILLER_265_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout692 _12560_/A vssd1 vssd1 vccd1 vccd1 _13655_/C1 sky130_fd_sc_hd__buf_4
X_13983_ _14033_/A1 _12978_/X _13982_/X _14037_/C1 vssd1 vssd1 vccd1 vccd1 _17956_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18510_ _19321_/CLK _18510_/D vssd1 vssd1 vccd1 vccd1 _18510_/Q sky130_fd_sc_hd__dfxtp_4
X_15722_ _15744_/A _15722_/B vssd1 vssd1 vccd1 vccd1 _15723_/B sky130_fd_sc_hd__and2_1
XFILLER_219_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12934_ _12933_/A _12822_/Y _12933_/Y vssd1 vssd1 vccd1 vccd1 _12934_/Y sky130_fd_sc_hd__a21oi_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _19490_/CLK _19490_/D vssd1 vssd1 vccd1 vccd1 _19490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15653_ _15653_/A _15653_/B vssd1 vssd1 vccd1 vccd1 _15653_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18441_ _19620_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _13978_/B vssd1 vssd1 vccd1 vccd1 _12865_/Y sky130_fd_sc_hd__inv_2
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _17696_/A0 _18411_/Q _14628_/S vssd1 vssd1 vccd1 vccd1 _18411_/D sky130_fd_sc_hd__mux2_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18372_ _19477_/CLK _18372_/D vssd1 vssd1 vccd1 vccd1 _18372_/Q sky130_fd_sc_hd__dfxtp_2
X_11816_ _11816_/A _12265_/B _09139_/X vssd1 vssd1 vccd1 vccd1 _11816_/X sky130_fd_sc_hd__or3b_4
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15584_ _15789_/A1 _15579_/Y _15580_/X _15789_/B1 vssd1 vssd1 vccd1 vccd1 _15584_/Y
+ sky130_fd_sc_hd__a31oi_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12796_ _12686_/X _12689_/X _12796_/S vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__mux2_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _19459_/Q _17377_/S vssd1 vssd1 vccd1 vccd1 _17323_/Y sky130_fd_sc_hd__nor2_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _18376_/Q _14559_/A2 _14559_/B1 input35/X vssd1 vssd1 vccd1 vccd1 _14536_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _18569_/Q _11759_/A2 _11909_/A _13125_/A vssd1 vssd1 vccd1 vccd1 _11747_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17254_ _19435_/Q _17256_/B _17253_/X vssd1 vssd1 vccd1 vccd1 _17255_/B sky130_fd_sc_hd__a21oi_1
X_14466_ _18318_/Q _17703_/A0 _14485_/S vssd1 vssd1 vccd1 vccd1 _18318_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11678_ _13411_/A _11678_/B vssd1 vssd1 vccd1 vccd1 _13443_/B sky130_fd_sc_hd__xnor2_4
XFILLER_105_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16205_ _16470_/A0 _18821_/Q _16225_/S vssd1 vssd1 vccd1 vccd1 _18821_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ _11293_/A _13316_/B _14156_/A0 vssd1 vssd1 vccd1 vccd1 _13417_/Y sky130_fd_sc_hd__a21oi_1
X_10629_ _10618_/S _10624_/X _10628_/X vssd1 vssd1 vccd1 vccd1 _10629_/X sky130_fd_sc_hd__o21a_1
X_17185_ _19413_/Q fanout536/X _17498_/A _17120_/B vssd1 vssd1 vccd1 vccd1 _17186_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_128_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14397_ _17704_/A0 _18248_/Q _14415_/S vssd1 vssd1 vccd1 vccd1 _18248_/D sky130_fd_sc_hd__mux2_1
X_16136_ _16142_/A1 _16135_/Y _16142_/B1 vssd1 vssd1 vccd1 vccd1 _18770_/D sky130_fd_sc_hd__a21oi_1
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13348_ _13791_/A _13346_/Y _13347_/X _13366_/B _13421_/A vssd1 vssd1 vccd1 vccd1
+ _13348_/X sky130_fd_sc_hd__a32o_1
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16067_ _16020_/A _16054_/A _16065_/Y _16066_/X _14427_/B vssd1 vssd1 vccd1 vccd1
+ _18739_/D sky130_fd_sc_hd__o221a_1
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13279_ _19435_/Q _12582_/X _13278_/X vssd1 vssd1 vccd1 vccd1 _13279_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15018_ _18507_/Q input207/X _16627_/S vssd1 vssd1 vccd1 vccd1 _18507_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16969_ _18773_/Q _16969_/A2 _16969_/B1 input239/X _16969_/C1 vssd1 vssd1 vccd1 vccd1
+ _16969_/X sky130_fd_sc_hd__a221o_1
XFILLER_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09510_ _09508_/X _09509_/X _10275_/S vssd1 vssd1 vccd1 vccd1 _09510_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18708_ _18761_/CLK _18708_/D vssd1 vssd1 vccd1 vccd1 _18708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09441_ _10264_/S _09440_/X _09439_/X _09463_/S vssd1 vssd1 vccd1 vccd1 _09441_/X
+ sky130_fd_sc_hd__a211o_1
X_18639_ _19142_/CLK _18639_/D vssd1 vssd1 vccd1 vccd1 _18639_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_213_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09372_ _18244_/Q _18819_/Q _09966_/S vssd1 vssd1 vccd1 vccd1 _09372_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput295 _11911_/X vssd1 vssd1 vccd1 vccd1 addr1[1] sky130_fd_sc_hd__buf_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09708_ _09708_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _09708_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10980_ _15526_/A vssd1 vssd1 vccd1 vccd1 _10980_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09639_ _09690_/A _09639_/B vssd1 vssd1 vccd1 vccd1 _09639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12650_ _10602_/A _12650_/B vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__and2b_1
XFILLER_231_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11601_ _11601_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11601_/Y sky130_fd_sc_hd__nand2_1
X_12581_ _12582_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _12581_/Y sky130_fd_sc_hd__nor2_8
XFILLER_70_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14320_ _18177_/Q _17704_/A0 _14338_/S vssd1 vssd1 vccd1 vccd1 _18177_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11532_ _13533_/A _11675_/B _11060_/Y vssd1 vssd1 vccd1 vccd1 _11674_/A sky130_fd_sc_hd__o21ai_4
XFILLER_278_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14251_ _18297_/Q _14261_/A2 _14250_/X _14449_/B vssd1 vssd1 vccd1 vccd1 _18123_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11463_ _11464_/C1 _11462_/X _11461_/X _09135_/S vssd1 vssd1 vccd1 vccd1 _11463_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202_ _13271_/C _13202_/B vssd1 vssd1 vccd1 vccd1 _13203_/A sky130_fd_sc_hd__or2_2
XFILLER_125_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10414_ _11333_/A1 _10414_/A2 _10413_/Y _11257_/C1 vssd1 vssd1 vccd1 vccd1 _10415_/B
+ sky130_fd_sc_hd__o211ai_4
X_14182_ _18702_/Q _18089_/Q _14200_/S vssd1 vssd1 vccd1 vccd1 _14183_/B sky130_fd_sc_hd__mux2_1
X_11394_ _19048_/Q _19016_/Q _11395_/C vssd1 vssd1 vccd1 vccd1 _11394_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13133_ _13135_/S _13131_/X _13132_/X _13129_/Y vssd1 vssd1 vccd1 vccd1 _13133_/X
+ sky130_fd_sc_hd__o22a_1
X_10345_ _18559_/Q _18434_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _10345_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18990_ _19118_/CLK _18990_/D vssd1 vssd1 vccd1 vccd1 _18990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _19496_/Q _13064_/B vssd1 vssd1 vccd1 vccd1 _13064_/X sky130_fd_sc_hd__or2_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _17951_/CLK _17941_/D vssd1 vssd1 vccd1 vccd1 _17941_/Q sky130_fd_sc_hd__dfxtp_4
X_10276_ _10294_/A1 _19582_/Q _10299_/S _19614_/Q _10300_/S vssd1 vssd1 vccd1 vccd1
+ _10276_/X sky130_fd_sc_hd__o221a_1
XFILLER_151_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1410 fanout1415/X vssd1 vssd1 vccd1 vccd1 _10099_/S sky130_fd_sc_hd__buf_6
X_12015_ _17782_/Q _17683_/A0 _12022_/S vssd1 vssd1 vccd1 vccd1 _17782_/D sky130_fd_sc_hd__mux2_1
XFILLER_266_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1421 _11403_/S vssd1 vssd1 vccd1 vccd1 _11477_/S sky130_fd_sc_hd__buf_6
Xfanout1432 _11484_/B1 vssd1 vssd1 vccd1 vccd1 _10180_/A sky130_fd_sc_hd__buf_8
X_17872_ _19324_/CLK _17872_/D vssd1 vssd1 vccd1 vccd1 _17872_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_266_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1443 _11002_/C1 vssd1 vssd1 vccd1 vccd1 _10335_/S sky130_fd_sc_hd__buf_8
Xfanout1454 _10337_/S1 vssd1 vssd1 vccd1 vccd1 _11001_/C1 sky130_fd_sc_hd__buf_6
XFILLER_227_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19611_ _19611_/CLK _19611_/D vssd1 vssd1 vccd1 vccd1 _19611_/Q sky130_fd_sc_hd__dfxtp_1
X_16823_ _17812_/Q _14672_/C _16836_/S vssd1 vssd1 vccd1 vccd1 _16981_/B sky130_fd_sc_hd__mux2_2
Xfanout1465 fanout1469/X vssd1 vssd1 vccd1 vccd1 _11340_/B2 sky130_fd_sc_hd__buf_6
XFILLER_266_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1476 _11125_/B2 vssd1 vssd1 vccd1 vccd1 _09797_/S sky130_fd_sc_hd__buf_6
Xfanout1487 _09885_/S vssd1 vssd1 vccd1 vccd1 _10054_/S sky130_fd_sc_hd__buf_6
XFILLER_285_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1498 _10290_/S vssd1 vssd1 vccd1 vccd1 _10281_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19542_ _19542_/CLK _19542_/D vssd1 vssd1 vccd1 vccd1 _19542_/Q sky130_fd_sc_hd__dfxtp_1
X_16754_ _19271_/Q _16754_/B vssd1 vssd1 vccd1 vccd1 _16759_/C sky130_fd_sc_hd__and2_2
X_13966_ _12442_/D _12752_/X _13965_/X _13966_/C1 vssd1 vssd1 vccd1 vccd1 _13966_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12917_ _15899_/A _12575_/Y _12909_/X _12916_/X vssd1 vssd1 vccd1 vccd1 _12917_/X
+ sky130_fd_sc_hd__a22o_1
X_15705_ _18588_/Q _15704_/C _18589_/Q vssd1 vssd1 vccd1 vccd1 _15706_/B sky130_fd_sc_hd__a21oi_1
X_16685_ _19248_/Q _16688_/C vssd1 vssd1 vccd1 vccd1 _16686_/B sky130_fd_sc_hd__and2_1
XFILLER_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19473_ _19507_/CLK _19473_/D vssd1 vssd1 vccd1 vccd1 _19473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13897_ _13895_/X _13896_/X _13893_/X vssd1 vssd1 vccd1 vccd1 _13897_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18424_ _19148_/CLK _18424_/D vssd1 vssd1 vccd1 vccd1 _18424_/Q sky130_fd_sc_hd__dfxtp_1
X_12848_ _17825_/Q _13942_/A2 _13942_/B1 _17857_/Q vssd1 vssd1 vccd1 vccd1 _12848_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15636_ _18125_/Q _15763_/A2 _15635_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _15687_/A
+ sky130_fd_sc_hd__o22a_2
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15567_ _19476_/Q _19410_/Q vssd1 vssd1 vccd1 vccd1 _15568_/B sky130_fd_sc_hd__or2_1
X_18355_ _19640_/CLK _18355_/D vssd1 vssd1 vccd1 vccd1 _18355_/Q sky130_fd_sc_hd__dfxtp_1
X_12779_ _15893_/A _12575_/Y _12778_/X vssd1 vssd1 vccd1 vccd1 _12779_/X sky130_fd_sc_hd__a21o_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _17720_/A0 _18368_/Q _14520_/S vssd1 vssd1 vccd1 vccd1 _18368_/D sky130_fd_sc_hd__mux2_1
XFILLER_147_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17306_ _17304_/Y _17305_/X _17210_/A vssd1 vssd1 vccd1 vccd1 _19452_/D sky130_fd_sc_hd__a21oi_1
XFILLER_222_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18286_ _19450_/CLK _18286_/D vssd1 vssd1 vccd1 vccd1 _18286_/Q sky130_fd_sc_hd__dfxtp_1
X_15498_ _19473_/Q _15497_/Y _15498_/S vssd1 vssd1 vccd1 vccd1 _15498_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17237_ _17235_/Y _17236_/X _17141_/A vssd1 vssd1 vccd1 vccd1 _19429_/D sky130_fd_sc_hd__a21oi_1
X_14449_ _18588_/Q _14449_/B vssd1 vssd1 vccd1 vccd1 _18301_/D sky130_fd_sc_hd__and2_1
XFILLER_174_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17168_ _17231_/A _17168_/B vssd1 vssd1 vccd1 vccd1 _19407_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16119_ _18762_/Q _16139_/B vssd1 vssd1 vccd1 vccd1 _16119_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09990_ input107/X input132/X _09990_/S vssd1 vssd1 vccd1 vccd1 _09991_/B sky130_fd_sc_hd__mux2_4
X_17099_ _19383_/Q _17115_/B vssd1 vssd1 vccd1 vccd1 _17099_/X sky130_fd_sc_hd__or2_1
XFILLER_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08941_ _17793_/Q _08941_/B vssd1 vssd1 vccd1 vccd1 _08941_/X sky130_fd_sc_hd__or2_2
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08872_ _17901_/Q _17899_/Q _08872_/C vssd1 vssd1 vccd1 vccd1 _12437_/A sky130_fd_sc_hd__or3_2
XFILLER_269_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_257_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09424_ _09424_/A _09424_/B vssd1 vssd1 vccd1 vccd1 _09424_/Y sky130_fd_sc_hd__nor2_1
XFILLER_240_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09355_ _19075_/Q _18979_/Q _11395_/C vssd1 vssd1 vccd1 vccd1 _09355_/X sky130_fd_sc_hd__mux2_1
XFILLER_240_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09286_ _18245_/Q _10217_/B _09285_/X _09374_/S vssd1 vssd1 vccd1 vccd1 _09286_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_179_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _18738_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_108_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _17865_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10130_ _19129_/Q _19161_/Q _10215_/S vssd1 vssd1 vccd1 vccd1 _10130_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10061_ _11365_/B2 _17659_/A0 _10060_/X _09523_/A vssd1 vssd1 vccd1 vccd1 _10061_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_134_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13820_ _19259_/Q _13943_/A2 _13943_/B1 _19291_/Q vssd1 vssd1 vccd1 vccd1 _13820_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13751_ _19449_/Q _13949_/A2 _13749_/X _13750_/X _13949_/C1 vssd1 vssd1 vccd1 vccd1
+ _13751_/X sky130_fd_sc_hd__o221a_1
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10963_ _10963_/A _10963_/B vssd1 vssd1 vccd1 vccd1 _10963_/Y sky130_fd_sc_hd__nor2_1
XFILLER_216_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ _12702_/A vssd1 vssd1 vccd1 vccd1 _12702_/Y sky130_fd_sc_hd__inv_2
X_16470_ _16470_/A0 _19077_/Q _16490_/S vssd1 vssd1 vccd1 vccd1 _19077_/D sky130_fd_sc_hd__mux2_1
XFILLER_203_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13682_ _17878_/Q _13747_/A2 _13681_/X _13682_/B2 vssd1 vssd1 vccd1 vccd1 _13682_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10894_ _18552_/Q _18427_/Q _18036_/Q _18004_/Q _11604_/S _11357_/S1 vssd1 vssd1
+ vccd1 vccd1 _10894_/X sky130_fd_sc_hd__mux4_1
XFILLER_203_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15421_ _15421_/A _15421_/B vssd1 vssd1 vccd1 vccd1 _15422_/B sky130_fd_sc_hd__xnor2_1
XPHY_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12633_ _12593_/A _12632_/X _12594_/X vssd1 vssd1 vccd1 vccd1 _12634_/B sky130_fd_sc_hd__o21a_1
XFILLER_71_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18140_ _18880_/CLK _18140_/D vssd1 vssd1 vccd1 vccd1 _18140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15352_ _18574_/Q _15388_/C vssd1 vssd1 vccd1 vccd1 _15352_/Y sky130_fd_sc_hd__nand2_1
X_12564_ _12584_/A _13167_/B vssd1 vssd1 vccd1 vccd1 _12564_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303_ _16621_/A0 _18162_/Q _14304_/S vssd1 vssd1 vccd1 vccd1 _18162_/D sky130_fd_sc_hd__mux2_1
X_11515_ _11428_/A _11514_/X _11515_/B1 vssd1 vssd1 vccd1 vccd1 _11515_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18071_ _19611_/CLK _18071_/D vssd1 vssd1 vccd1 vccd1 _18071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15283_ _18570_/Q _15351_/A2 _15282_/X _17338_/A vssd1 vssd1 vccd1 vccd1 _18570_/D
+ sky130_fd_sc_hd__o211a_1
X_12495_ _12578_/A _12544_/A vssd1 vssd1 vccd1 vccd1 _12495_/Y sky130_fd_sc_hd__nor2_4
XFILLER_138_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17022_ _17178_/B _17046_/A2 _17021_/X _17354_/A vssd1 vssd1 vccd1 vccd1 _19347_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14234_ _18115_/Q _14260_/B vssd1 vssd1 vccd1 vccd1 _14234_/X sky130_fd_sc_hd__or2_1
XFILLER_8_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11446_ _13357_/S _11446_/B vssd1 vssd1 vccd1 vccd1 _13351_/A sky130_fd_sc_hd__nor2_8
XFILLER_172_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14165_ _18774_/Q _16141_/B _16145_/B vssd1 vssd1 vccd1 vccd1 _14204_/S sky130_fd_sc_hd__or3_4
XFILLER_166_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11377_ _18984_/Q _11479_/B vssd1 vssd1 vccd1 vccd1 _11377_/X sky130_fd_sc_hd__or2_1
XFILLER_166_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13116_ _13116_/A _13116_/B vssd1 vssd1 vccd1 vccd1 _13116_/Y sky130_fd_sc_hd__nor2_1
XFILLER_180_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10328_ _10334_/A1 _19581_/Q _09179_/B _19613_/Q vssd1 vssd1 vccd1 vccd1 _10328_/X
+ sky130_fd_sc_hd__o22a_1
X_14096_ _16314_/A0 _18036_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _18036_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18973_ _18973_/CLK _18973_/D vssd1 vssd1 vccd1 vccd1 _18973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17924_ _17930_/CLK _17924_/D vssd1 vssd1 vccd1 vccd1 _17924_/Q sky130_fd_sc_hd__dfxtp_4
X_13047_ _13047_/A vssd1 vssd1 vccd1 vccd1 _13047_/Y sky130_fd_sc_hd__inv_2
X_10259_ _10257_/X _10258_/X _10264_/S vssd1 vssd1 vccd1 vccd1 _10259_/X sky130_fd_sc_hd__mux2_1
XFILLER_252_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1240 _09108_/X vssd1 vssd1 vccd1 vccd1 _11257_/C1 sky130_fd_sc_hd__buf_12
Xfanout1251 _10905_/S vssd1 vssd1 vccd1 vccd1 _13739_/A sky130_fd_sc_hd__buf_12
XFILLER_266_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17855_ _19268_/CLK _17855_/D vssd1 vssd1 vccd1 vccd1 _17855_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1262 _13807_/A vssd1 vssd1 vccd1 vccd1 _13237_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout1273 _12276_/X vssd1 vssd1 vccd1 vccd1 _12277_/B sky130_fd_sc_hd__buf_6
XFILLER_94_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1284 _16002_/A2 vssd1 vssd1 vccd1 vccd1 _15918_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_226_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16806_ _19290_/Q _16807_/C _19291_/Q vssd1 vssd1 vccd1 vccd1 _16808_/B sky130_fd_sc_hd__a21oi_1
Xfanout1295 _14586_/A vssd1 vssd1 vccd1 vccd1 _14596_/A sky130_fd_sc_hd__buf_4
XFILLER_226_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17786_ _19159_/CLK _17786_/D vssd1 vssd1 vccd1 vccd1 _17786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14998_ _14998_/A vssd1 vssd1 vccd1 vccd1 _14998_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_35_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19525_ _19525_/CLK _19525_/D vssd1 vssd1 vccd1 vccd1 _19525_/Q sky130_fd_sc_hd__dfxtp_1
X_16737_ _16737_/A _16743_/C vssd1 vssd1 vccd1 vccd1 _16737_/Y sky130_fd_sc_hd__nor2_1
XFILLER_223_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13949_ _19455_/Q _13949_/A2 _13947_/X _13948_/X _13949_/C1 vssd1 vssd1 vccd1 vccd1
+ _13949_/X sky130_fd_sc_hd__o221a_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19456_ _19458_/CLK _19456_/D vssd1 vssd1 vccd1 vccd1 _19456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16668_ _16768_/A _16674_/C vssd1 vssd1 vccd1 vccd1 _16668_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18407_ _19197_/CLK _18407_/D vssd1 vssd1 vccd1 vccd1 _18407_/Q sky130_fd_sc_hd__dfxtp_1
X_15619_ _15620_/A _15620_/B _15638_/D vssd1 vssd1 vccd1 vccd1 _15619_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19387_ _19546_/CLK _19387_/D vssd1 vssd1 vccd1 vccd1 _19387_/Q sky130_fd_sc_hd__dfxtp_1
X_16599_ _17699_/A0 _19202_/Q _16622_/S vssd1 vssd1 vccd1 vccd1 _19202_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09140_ _15549_/A _09139_/X _09140_/S vssd1 vssd1 vccd1 vccd1 _09144_/C sky130_fd_sc_hd__mux2_1
X_18338_ _19618_/CLK _18338_/D vssd1 vssd1 vccd1 vccd1 _18338_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_6_wb_clk_i _19652_/A vssd1 vssd1 vccd1 vccd1 _19118_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_175_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09071_ _17901_/Q _12264_/B vssd1 vssd1 vccd1 vccd1 _12455_/A sky130_fd_sc_hd__nor2_4
X_18269_ _18272_/CLK _18269_/D vssd1 vssd1 vccd1 vccd1 _18269_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_201_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19639_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_190_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09973_ _19068_/Q _18972_/Q _09973_/S vssd1 vssd1 vccd1 vccd1 _09973_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08924_ _16525_/A _14074_/C _14074_/B vssd1 vssd1 vccd1 vccd1 _11985_/C sky130_fd_sc_hd__and3_2
XFILLER_131_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08855_ _17795_/Q vssd1 vssd1 vccd1 vccd1 _14741_/A sky130_fd_sc_hd__inv_2
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09407_ _10294_/A1 _19593_/Q _19561_/Q _09428_/B2 vssd1 vssd1 vccd1 vccd1 _09407_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09338_ _18540_/Q _18415_/Q _09344_/S vssd1 vssd1 vccd1 vccd1 _09338_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09269_ _19076_/Q _18980_/Q _09269_/S vssd1 vssd1 vccd1 vccd1 _09269_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11300_ _18985_/Q _11300_/B vssd1 vssd1 vccd1 vccd1 _11300_/X sky130_fd_sc_hd__or2_1
XFILLER_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12280_ _18092_/Q _12305_/A2 _14692_/A2 _18515_/Q vssd1 vssd1 vccd1 vccd1 _12476_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_181_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11231_ _18547_/Q _11247_/S vssd1 vssd1 vccd1 vccd1 _11231_/X sky130_fd_sc_hd__or2_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11162_ _19051_/Q _19019_/Q _11171_/S vssd1 vssd1 vccd1 vccd1 _11162_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _11017_/A1 _19161_/Q _10176_/S _19129_/Q vssd1 vssd1 vccd1 vccd1 _10113_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ _18700_/Q _15970_/A2 _15976_/B1 _18749_/Q _15976_/C1 vssd1 vssd1 vccd1 vccd1
+ _15970_/X sky130_fd_sc_hd__a221o_1
X_11093_ _10930_/S _11092_/X _11583_/A vssd1 vssd1 vccd1 vccd1 _11093_/X sky130_fd_sc_hd__a21o_1
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10044_ _15481_/A _10037_/X _11286_/B1 vssd1 vssd1 vccd1 vccd1 _10044_/Y sky130_fd_sc_hd__a21oi_1
X_14921_ _17813_/Q _15002_/B vssd1 vssd1 vccd1 vccd1 _14921_/X sky130_fd_sc_hd__or2_1
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_wb_clk_i clkbuf_leaf_78_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19627_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17640_ _17706_/A0 _19568_/Q _17657_/S vssd1 vssd1 vccd1 vccd1 _19568_/D sky130_fd_sc_hd__mux2_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14852_ _19229_/Q _15014_/B _14934_/C _14934_/D vssd1 vssd1 vccd1 vccd1 _14852_/X
+ sky130_fd_sc_hd__and4_4
XFILLER_236_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13803_ _18126_/Q _13802_/C _18127_/Q vssd1 vssd1 vccd1 vccd1 _13804_/B sky130_fd_sc_hd__a21oi_1
X_17571_ _17571_/A _17583_/B vssd1 vssd1 vccd1 vccd1 _17571_/X sky130_fd_sc_hd__or2_1
X_14783_ _14875_/A1 _14782_/X _14865_/B1 vssd1 vssd1 vccd1 vccd1 _14783_/Y sky130_fd_sc_hd__o21ai_2
X_11995_ _17762_/Q _17663_/A0 _12019_/S vssd1 vssd1 vccd1 vccd1 _17762_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19310_ _19310_/CLK _19310_/D vssd1 vssd1 vccd1 vccd1 _19310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16522_ _16522_/A0 _19128_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _19128_/D sky130_fd_sc_hd__mux2_1
X_13734_ _13968_/A1 _13726_/X _13733_/X _13323_/B vssd1 vssd1 vccd1 vccd1 _13734_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10946_ _09107_/D _10935_/X _10943_/X _10945_/X vssd1 vssd1 vccd1 vccd1 _10946_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_204_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19241_ _19280_/CLK _19241_/D vssd1 vssd1 vccd1 vccd1 _19241_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16453_ _19061_/Q _16618_/A0 _16453_/S vssd1 vssd1 vccd1 vccd1 _19061_/D sky130_fd_sc_hd__mux2_1
X_13665_ _13665_/A _13665_/B vssd1 vssd1 vccd1 vccd1 _14149_/B sky130_fd_sc_hd__xnor2_2
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10877_ _11596_/A1 _19638_/Q _18927_/Q _11604_/S vssd1 vssd1 vccd1 vccd1 _10877_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15404_/A _15404_/B vssd1 vssd1 vccd1 vccd1 _15404_/Y sky130_fd_sc_hd__nor2_1
X_12616_ _11739_/A _12610_/B _13083_/B vssd1 vssd1 vccd1 vccd1 _12616_/X sky130_fd_sc_hd__o21a_1
X_19172_ _19627_/CLK _19172_/D vssd1 vssd1 vccd1 vccd1 _19172_/Q sky130_fd_sc_hd__dfxtp_1
X_16384_ _10532_/B _18995_/Q _16391_/S vssd1 vssd1 vccd1 vccd1 _18995_/D sky130_fd_sc_hd__mux2_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13758_/A _13581_/X _13956_/B1 vssd1 vssd1 vccd1 vccd1 _13596_/X sky130_fd_sc_hd__a21o_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18123_ _19450_/CLK _18123_/D vssd1 vssd1 vccd1 vccd1 _18123_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15335_ _15336_/B _15335_/B vssd1 vssd1 vccd1 vccd1 _15335_/X sky130_fd_sc_hd__and2b_1
X_12547_ _17855_/Q _12919_/A2 _12546_/X _13945_/B2 _13115_/C1 vssd1 vssd1 vccd1 vccd1
+ _12547_/X sky130_fd_sc_hd__a221o_1
XFILLER_184_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18054_ _18632_/CLK _18054_/D vssd1 vssd1 vccd1 vccd1 _18054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15266_ _15171_/A _15171_/B _15263_/X _15265_/X vssd1 vssd1 vccd1 vccd1 _15268_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_117_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12478_ _12483_/A _12478_/B vssd1 vssd1 vccd1 vccd1 _12478_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_3 _18198_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17005_ _19339_/Q _17009_/B vssd1 vssd1 vccd1 vccd1 _17005_/X sky130_fd_sc_hd__or2_1
X_14217_ _18280_/Q _14252_/B _14216_/X _16046_/A vssd1 vssd1 vccd1 vccd1 _18106_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11429_ _18639_/Q _18061_/Q _19080_/Q _18984_/Q _11503_/S0 _11503_/S1 vssd1 vssd1
+ vccd1 vccd1 _11429_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15197_ _17913_/Q _15369_/A vssd1 vssd1 vccd1 vccd1 _15199_/B sky130_fd_sc_hd__and2_1
X_14148_ _14148_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14149_/D sky130_fd_sc_hd__or2_1
XFILLER_259_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18956_ _19118_/CLK _18956_/D vssd1 vssd1 vccd1 vccd1 _18956_/Q sky130_fd_sc_hd__dfxtp_1
X_14079_ _16595_/A0 _18019_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _18019_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17907_ _18881_/CLK _17907_/D vssd1 vssd1 vccd1 vccd1 _17907_/Q sky130_fd_sc_hd__dfxtp_4
X_18887_ _19208_/CLK _18887_/D vssd1 vssd1 vccd1 vccd1 _18887_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1070 _14027_/A2 vssd1 vssd1 vccd1 vccd1 _14036_/A sky130_fd_sc_hd__buf_4
XFILLER_94_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1081 _09980_/A2 vssd1 vssd1 vccd1 vccd1 _16461_/A0 sky130_fd_sc_hd__clkbuf_2
X_17838_ _19310_/CLK _17838_/D vssd1 vssd1 vccd1 vccd1 _17838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1092 _09743_/B vssd1 vssd1 vccd1 vccd1 _16529_/A0 sky130_fd_sc_hd__buf_2
XFILLER_254_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17769_ _19565_/CLK _17769_/D vssd1 vssd1 vccd1 vccd1 _17769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19508_ _19521_/CLK _19508_/D vssd1 vssd1 vccd1 vccd1 _19508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19439_ _19543_/CLK _19439_/D vssd1 vssd1 vccd1 vccd1 _19439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09123_ _09129_/S _09121_/X _09122_/X _12408_/A vssd1 vssd1 vccd1 vccd1 _09123_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09054_ _09053_/Y _09052_/Y _08945_/X _17931_/Q vssd1 vssd1 vccd1 vccd1 _09054_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_163_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09956_ _11190_/A1 _18134_/Q _18780_/Q _09973_/S vssd1 vssd1 vccd1 vccd1 _09956_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08907_ _08932_/A _12053_/A _17802_/Q _12051_/A vssd1 vssd1 vccd1 vccd1 _08907_/Y
+ sky130_fd_sc_hd__o31ai_2
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _19069_/Q _18973_/Q _10496_/B vssd1 vssd1 vccd1 vccd1 _09887_/X sky130_fd_sc_hd__mux2_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _09031_/S vssd1 vssd1 vccd1 vccd1 _09028_/B sky130_fd_sc_hd__clkinv_4
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_404 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_415 _13647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_426 _11822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10800_ _18647_/Q _11605_/S vssd1 vssd1 vccd1 vccd1 _10800_/X sky130_fd_sc_hd__or2_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_437 _13019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_448 _13637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11780_ _11869_/B _11859_/B _11774_/B _11779_/X vssd1 vssd1 vccd1 vccd1 _11780_/X
+ sky130_fd_sc_hd__o211a_4
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_459 _18646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10731_ _11622_/C1 _10725_/X _10728_/X _10730_/X _11508_/B1 vssd1 vssd1 vccd1 vccd1
+ _10731_/X sky130_fd_sc_hd__a311o_2
XFILLER_41_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_194_wb_clk_i clkbuf_4_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19644_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13450_ _17871_/Q _13747_/A2 _13448_/X _13747_/B2 vssd1 vssd1 vccd1 vccd1 _13450_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10662_ _10662_/A1 _18156_/Q _18802_/Q _10667_/S vssd1 vssd1 vccd1 vccd1 _10662_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _09457_/B _12412_/A _12400_/Y _14001_/C1 vssd1 vssd1 vccd1 vccd1 _17908_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_123_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19323_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13381_ _13920_/B2 _13370_/X _13380_/X vssd1 vssd1 vccd1 vccd1 _14002_/B sky130_fd_sc_hd__a21oi_4
XFILLER_210_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10593_ _10591_/X _10592_/X _10668_/S vssd1 vssd1 vccd1 vccd1 _10594_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15120_ _15120_/A _15120_/B vssd1 vssd1 vccd1 vccd1 _15120_/Y sky130_fd_sc_hd__nor2_2
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12332_ _17803_/Q _17802_/Q _17801_/Q _12332_/D vssd1 vssd1 vccd1 vccd1 _12333_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _18535_/Q _17662_/A0 _15079_/S vssd1 vssd1 vccd1 vccd1 _18535_/D sky130_fd_sc_hd__mux2_1
X_12263_ _12263_/A vssd1 vssd1 vccd1 vccd1 _15328_/B sky130_fd_sc_hd__inv_2
XFILLER_181_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14002_ _14028_/A _14002_/B vssd1 vssd1 vccd1 vccd1 _14002_/Y sky130_fd_sc_hd__nand2_1
X_11214_ _11214_/A _11214_/B vssd1 vssd1 vccd1 vccd1 _11215_/B sky130_fd_sc_hd__nor2_4
X_12194_ _17862_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12200_/C sky130_fd_sc_hd__and2_2
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18810_ _19607_/CLK _18810_/D vssd1 vssd1 vccd1 vccd1 _18810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11145_ _18987_/Q _11224_/B vssd1 vssd1 vccd1 vccd1 _11145_/X sky130_fd_sc_hd__or2_1
XFILLER_68_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18741_ _18741_/CLK _18741_/D vssd1 vssd1 vccd1 vccd1 _18741_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_283_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15953_ _15953_/A _15953_/B vssd1 vssd1 vccd1 vccd1 _15953_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11076_ _18424_/Q _11300_/B _11075_/X _11562_/S vssd1 vssd1 vccd1 vccd1 _11076_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput140 dout1[3] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput151 dout1[4] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_hd__clkbuf_2
XFILLER_264_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput162 dout1[5] vssd1 vssd1 vccd1 vccd1 input162/X sky130_fd_sc_hd__clkbuf_2
X_10027_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10027_/Y sky130_fd_sc_hd__nand2_1
X_14904_ _18122_/Q _14893_/S _14852_/X _14903_/X vssd1 vssd1 vccd1 vccd1 _14904_/X
+ sky130_fd_sc_hd__o211a_2
X_18672_ _18683_/CLK _18672_/D vssd1 vssd1 vccd1 vccd1 _18672_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput173 irq[11] vssd1 vssd1 vccd1 vccd1 _15088_/C sky130_fd_sc_hd__clkbuf_2
X_15884_ _15884_/A _15905_/B _15908_/C vssd1 vssd1 vccd1 vccd1 _15884_/X sky130_fd_sc_hd__and3_1
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput184 irq[7] vssd1 vssd1 vccd1 vccd1 _15085_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 localMemory_wb_adr_i[14] vssd1 vssd1 vccd1 vccd1 input195/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17623_ _19391_/Q _15092_/B input177/X _17592_/X _17623_/B1 vssd1 vssd1 vccd1 vccd1
+ _17623_/X sky130_fd_sc_hd__a41o_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _14835_/A vssd1 vssd1 vccd1 vccd1 _14835_/Y sky130_fd_sc_hd__inv_2
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _19521_/Q _17493_/B _17553_/X vssd1 vssd1 vccd1 vccd1 _19521_/D sky130_fd_sc_hd__o21ba_1
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14766_ _14763_/Y _14765_/Y _14879_/B1 vssd1 vssd1 vccd1 vccd1 _14766_/Y sky130_fd_sc_hd__a21oi_4
X_11978_ _18736_/Q _18735_/Q _18733_/Q vssd1 vssd1 vccd1 vccd1 _11979_/C sky130_fd_sc_hd__or3b_2
XFILLER_147_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ _16538_/A0 _19111_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _19111_/D sky130_fd_sc_hd__mux2_1
XFILLER_220_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10929_ _19637_/Q _18926_/Q _10929_/S vssd1 vssd1 vccd1 vccd1 _10929_/X sky130_fd_sc_hd__mux2_1
X_13717_ _19514_/Q _13947_/A2 _13781_/B1 _13716_/X vssd1 vssd1 vccd1 vccd1 _13717_/X
+ sky130_fd_sc_hd__o211a_1
X_17485_ _13566_/A _17520_/A2 _17532_/A2 _17809_/Q _17550_/A vssd1 vssd1 vccd1 vccd1
+ _17485_/X sky130_fd_sc_hd__a221o_1
X_14697_ input43/X input68/X _14784_/S vssd1 vssd1 vccd1 vccd1 _14698_/B sky130_fd_sc_hd__mux2_8
XFILLER_32_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19224_ _19647_/CLK _19224_/D vssd1 vssd1 vccd1 vccd1 _19224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16436_ _19044_/Q _17668_/A0 _16457_/S vssd1 vssd1 vccd1 vccd1 _19044_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13648_ _17845_/Q _13744_/A2 _13744_/B1 _17877_/Q vssd1 vssd1 vccd1 vccd1 _13648_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19155_/CLK _19155_/D vssd1 vssd1 vccd1 vccd1 _19155_/Q sky130_fd_sc_hd__dfxtp_1
X_16367_ _16500_/A0 _18978_/Q _16388_/S vssd1 vssd1 vccd1 vccd1 _18978_/D sky130_fd_sc_hd__mux2_1
X_13579_ _13579_/A _13579_/B _13577_/X vssd1 vssd1 vccd1 vccd1 _13579_/X sky130_fd_sc_hd__or3b_4
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18106_ _18734_/CLK _18106_/D vssd1 vssd1 vccd1 vccd1 _18106_/Q sky130_fd_sc_hd__dfxtp_4
X_15318_ _15369_/A _15313_/Y _15317_/Y vssd1 vssd1 vccd1 vccd1 _15318_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_258_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16298_ _17696_/A0 _18911_/Q _16323_/S vssd1 vssd1 vccd1 vccd1 _18911_/D sky130_fd_sc_hd__mux2_1
X_19086_ _19118_/CLK _19086_/D vssd1 vssd1 vccd1 vccd1 _19086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18037_ _19600_/CLK _18037_/D vssd1 vssd1 vccd1 vccd1 _18037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15249_ _12788_/B _15248_/Y _15307_/B vssd1 vssd1 vccd1 vccd1 _15250_/C sky130_fd_sc_hd__a21oi_2
XFILLER_160_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09810_ _11622_/A1 _09799_/X _09809_/X _11621_/C1 vssd1 vssd1 vccd1 vccd1 _09810_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09741_ _10085_/A _09047_/X _09737_/X _09740_/X vssd1 vssd1 vccd1 vccd1 _09741_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_140_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18939_ _19099_/CLK _18939_/D vssd1 vssd1 vccd1 vccd1 _18939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_268_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09672_ _11172_/A1 _19199_/Q _19167_/Q _09688_/S _11480_/C1 vssd1 vssd1 vccd1 vccd1
+ _09672_/X sky130_fd_sc_hd__a221o_1
XFILLER_283_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09106_ _10632_/S _09106_/B vssd1 vssd1 vccd1 vccd1 _09108_/D sky130_fd_sc_hd__nand2_1
XFILLER_202_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09037_ _09034_/B _09036_/X _09326_/A vssd1 vssd1 vccd1 vccd1 _09037_/X sky130_fd_sc_hd__a21o_1
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1806 _14442_/B vssd1 vssd1 vccd1 vccd1 _14452_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_278_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1817 _17366_/A vssd1 vssd1 vccd1 vccd1 _17106_/C1 sky130_fd_sc_hd__buf_2
XFILLER_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout830 _16476_/A0 vssd1 vssd1 vccd1 vccd1 _17708_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout1828 _17336_/A vssd1 vssd1 vccd1 vccd1 _17360_/A sky130_fd_sc_hd__buf_4
Xfanout841 _10989_/X vssd1 vssd1 vccd1 vccd1 _16610_/A0 sky130_fd_sc_hd__clkbuf_8
Xfanout1839 _14179_/A vssd1 vssd1 vccd1 vccd1 _14177_/A sky130_fd_sc_hd__buf_4
XFILLER_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout852 _10792_/A2 vssd1 vssd1 vccd1 vccd1 _17680_/A0 sky130_fd_sc_hd__clkbuf_4
X_09939_ _08843_/A _09927_/X _09938_/X _10264_/S _10996_/B1 vssd1 vssd1 vccd1 vccd1
+ _09939_/X sky130_fd_sc_hd__o221a_1
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout863 _10609_/X vssd1 vssd1 vccd1 vccd1 _16549_/A0 sky130_fd_sc_hd__clkbuf_2
Xfanout874 _17721_/A0 vssd1 vssd1 vccd1 vccd1 _17688_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout885 _10028_/X vssd1 vssd1 vccd1 vccd1 _12796_/S sky130_fd_sc_hd__buf_4
Xfanout896 _16203_/A0 vssd1 vssd1 vccd1 vccd1 _17700_/A0 sky130_fd_sc_hd__clkbuf_4
X_12950_ _12936_/S _12710_/X _12746_/X vssd1 vssd1 vccd1 vccd1 _12990_/B sky130_fd_sc_hd__o21ai_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11901_ _11901_/A _11901_/B vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__or2_1
XFILLER_100_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _12705_/X _12713_/X _12935_/S vssd1 vssd1 vccd1 vccd1 _12881_/X sky130_fd_sc_hd__mux2_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_201 _14036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _17906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 _18383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _16314_/A0 _18427_/Q _14631_/S vssd1 vssd1 vccd1 vccd1 _18427_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11832_ _11832_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__nor2_2
XANTENNA_234 _18392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 _18725_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_256 _15854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_267 input226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _18384_/Q _14575_/A2 _14575_/B1 input12/X vssd1 vssd1 vccd1 vccd1 _14552_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_278 input243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _18581_/Q _14349_/B _11769_/B1 _13566_/A vssd1 vssd1 vccd1 vccd1 _11763_/X
+ sky130_fd_sc_hd__a22o_4
XANTENNA_289 _11931_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _19377_/Q _13951_/A2 _13500_/X _13501_/X _13951_/C1 vssd1 vssd1 vccd1 vccd1
+ _13502_/X sky130_fd_sc_hd__o221a_4
X_10714_ _11024_/A1 _10712_/X _10713_/X vssd1 vssd1 vccd1 vccd1 _11864_/A sky130_fd_sc_hd__o21ai_4
X_14482_ _18334_/Q _17686_/A0 _14485_/S vssd1 vssd1 vccd1 vccd1 _18334_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _17268_/Y _17269_/X _17285_/A vssd1 vssd1 vccd1 vccd1 _19440_/D sky130_fd_sc_hd__a21oi_1
X_11694_ _12432_/B1 _14525_/A vssd1 vssd1 vccd1 vccd1 _11694_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16221_ _17718_/A0 _18837_/Q _16226_/S vssd1 vssd1 vccd1 vccd1 _18837_/D sky130_fd_sc_hd__mux2_1
X_13433_ _19375_/Q _13951_/A2 _13431_/X _13432_/X _13951_/C1 vssd1 vssd1 vccd1 vccd1
+ _13433_/X sky130_fd_sc_hd__o221a_4
X_10645_ _18039_/Q _18007_/Q _10645_/S vssd1 vssd1 vccd1 vccd1 _10645_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16152_ _18775_/Q _16146_/X _16151_/X vssd1 vssd1 vccd1 vccd1 _18775_/D sky130_fd_sc_hd__o21ba_1
XFILLER_167_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13364_ _15429_/A2 _13361_/X _13363_/A _13936_/B2 vssd1 vssd1 vccd1 vccd1 _13365_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10576_ _10662_/A1 _18228_/Q _10650_/S _18963_/Q _10649_/A1 vssd1 vssd1 vccd1 vccd1
+ _10576_/X sky130_fd_sc_hd__o221a_1
XFILLER_154_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15103_ _18778_/Q _18777_/Q vssd1 vssd1 vccd1 vccd1 _15103_/Y sky130_fd_sc_hd__nor2_4
X_12315_ _12439_/A _12315_/B vssd1 vssd1 vccd1 vccd1 _13260_/B sky130_fd_sc_hd__or2_4
X_16083_ _18744_/Q _16093_/B vssd1 vssd1 vccd1 vccd1 _16083_/Y sky130_fd_sc_hd__nand2_1
XFILLER_182_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13295_ _15357_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _13295_/Y sky130_fd_sc_hd__nand2_1
X_15034_ _18523_/Q input200/X _15038_/S vssd1 vssd1 vccd1 vccd1 _18523_/D sky130_fd_sc_hd__mux2_1
XFILLER_182_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12246_ _17881_/Q _12248_/C _12245_/Y vssd1 vssd1 vccd1 vccd1 _17881_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_91_wb_clk_i clkbuf_leaf_91_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _18746_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12177_ _12203_/A _12177_/B _12178_/B vssd1 vssd1 vccd1 vccd1 _17855_/D sky130_fd_sc_hd__nor3_1
XFILLER_174_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_wb_clk_i clkbuf_4_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19618_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11128_ _10040_/S _11127_/X _11623_/A1 vssd1 vssd1 vccd1 vccd1 _11128_/X sky130_fd_sc_hd__a21o_1
XFILLER_268_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16985_ _19329_/Q _17043_/B vssd1 vssd1 vccd1 vccd1 _16985_/X sky130_fd_sc_hd__or2_1
XFILLER_49_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18724_ _18775_/CLK _18724_/D vssd1 vssd1 vccd1 vccd1 _18724_/Q sky130_fd_sc_hd__dfxtp_1
X_15936_ _18687_/Q _15948_/A2 _15948_/B1 _15935_/X _15945_/C1 vssd1 vssd1 vccd1 vccd1
+ _15936_/X sky130_fd_sc_hd__a221o_1
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ _12594_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _13535_/S sky130_fd_sc_hd__and2_4
XFILLER_260_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18655_ _19076_/CLK _18655_/D vssd1 vssd1 vccd1 vccd1 _18655_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15867_ _18664_/Q _15853_/Y _15906_/B1 vssd1 vssd1 vccd1 vccd1 _15867_/X sky130_fd_sc_hd__a21o_1
XFILLER_236_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17606_ _19544_/Q _17624_/A2 _17591_/X _17187_/B _17605_/X vssd1 vssd1 vccd1 vccd1
+ _19544_/D sky130_fd_sc_hd__o221a_1
X_14818_ _18483_/Q _15001_/A2 _14817_/Y _12249_/A vssd1 vssd1 vccd1 vccd1 _18483_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18586_ _19448_/CLK _18586_/D vssd1 vssd1 vccd1 vccd1 _18586_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ _19487_/Q _15781_/S _15796_/Y _17208_/A vssd1 vssd1 vccd1 vccd1 _15798_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17537_ _17819_/Q _17543_/B1 _17531_/B _13904_/B vssd1 vssd1 vccd1 vccd1 _17538_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14749_ _18476_/Q _14720_/A _14748_/Y _12241_/A vssd1 vssd1 vccd1 vccd1 _18476_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17468_ _17468_/A _17547_/B vssd1 vssd1 vccd1 vccd1 _17468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19207_ _19587_/CLK _19207_/D vssd1 vssd1 vccd1 vccd1 _19207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16419_ _16617_/A0 _19028_/Q _16420_/S vssd1 vssd1 vccd1 vccd1 _19028_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17399_ _17123_/Y _17462_/B _17398_/Y _17141_/A vssd1 vssd1 vccd1 vccd1 _17399_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_285_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19138_ _19138_/CLK _19138_/D vssd1 vssd1 vccd1 vccd1 _19138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19069_ _19588_/CLK _19069_/D vssd1 vssd1 vccd1 vccd1 _19069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput400 _11951_/X vssd1 vssd1 vccd1 vccd1 din0[31] sky130_fd_sc_hd__buf_4
Xoutput411 _18481_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[10] sky130_fd_sc_hd__buf_4
Xoutput422 _18491_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[20] sky130_fd_sc_hd__buf_4
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput433 _18501_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[30] sky130_fd_sc_hd__buf_4
Xoutput444 _08881_/X vssd1 vssd1 vccd1 vccd1 probe_env[1] sky130_fd_sc_hd__buf_4
Xoutput455 _18115_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[14] sky130_fd_sc_hd__buf_4
XFILLER_114_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput466 _18125_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[24] sky130_fd_sc_hd__buf_4
XFILLER_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput477 _18106_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[5] sky130_fd_sc_hd__buf_4
XFILLER_99_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09724_ _19071_/Q _18975_/Q _09724_/S vssd1 vssd1 vccd1 vccd1 _09724_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09655_ input127/X input163/X _09655_/S vssd1 vssd1 vccd1 vccd1 _09655_/X sky130_fd_sc_hd__mux2_8
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09586_ _10742_/A1 _09582_/X _09583_/X vssd1 vssd1 vccd1 vccd1 _09586_/X sky130_fd_sc_hd__o21a_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10430_ _11510_/S1 _10419_/X _10429_/X _11438_/B1 vssd1 vssd1 vccd1 vccd1 _10430_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10361_ _18263_/Q _18838_/Q _10370_/S vssd1 vssd1 vccd1 vccd1 _10361_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12100_ _17826_/Q _17827_/Q _12100_/C vssd1 vssd1 vccd1 vccd1 _12106_/C sky130_fd_sc_hd__and3_2
XFILLER_136_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13080_ _13254_/B2 _13081_/A _13057_/Y _13079_/X vssd1 vssd1 vccd1 vccd1 _13080_/X
+ sky130_fd_sc_hd__a211o_1
X_10292_ _18903_/Q _10364_/B vssd1 vssd1 vccd1 vccd1 _10292_/X sky130_fd_sc_hd__or2_1
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12031_ _17793_/Q _12073_/B vssd1 vssd1 vccd1 vccd1 _12031_/X sky130_fd_sc_hd__or2_1
XFILLER_104_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1603 _17550_/A vssd1 vssd1 vccd1 vccd1 _17538_/A sky130_fd_sc_hd__buf_4
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1614 _11711_/A vssd1 vssd1 vccd1 vccd1 _15014_/B sky130_fd_sc_hd__buf_6
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1625 _09650_/B1 vssd1 vssd1 vccd1 vccd1 _11692_/A1 sky130_fd_sc_hd__buf_4
Xfanout1636 _12420_/A1 vssd1 vssd1 vccd1 vccd1 _12429_/A1 sky130_fd_sc_hd__buf_12
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1647 _11618_/A1 vssd1 vssd1 vccd1 vccd1 _11284_/A1 sky130_fd_sc_hd__buf_6
XFILLER_266_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1658 _11506_/A1 vssd1 vssd1 vccd1 vccd1 _11512_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_238_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout660 _12569_/Y vssd1 vssd1 vccd1 vccd1 _13243_/B1 sky130_fd_sc_hd__buf_6
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout671 _11649_/Y vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__buf_4
XFILLER_247_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1669 _09958_/C1 vssd1 vssd1 vccd1 vccd1 _15481_/A sky130_fd_sc_hd__clkbuf_16
X_16770_ _19277_/Q _16770_/B vssd1 vssd1 vccd1 vccd1 _16775_/C sky130_fd_sc_hd__and2_2
Xfanout682 _13950_/C1 vssd1 vssd1 vccd1 vccd1 _13883_/C1 sky130_fd_sc_hd__buf_6
X_13982_ _17956_/Q _14020_/B vssd1 vssd1 vccd1 vccd1 _13982_/X sky130_fd_sc_hd__or2_1
Xfanout693 _12557_/X vssd1 vssd1 vccd1 vccd1 _12560_/A sky130_fd_sc_hd__buf_6
XFILLER_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15721_ _15744_/A _15722_/B vssd1 vssd1 vccd1 vccd1 _15723_/A sky130_fd_sc_hd__nor2_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12933_ _12933_/A _12933_/B vssd1 vssd1 vccd1 vccd1 _12933_/Y sky130_fd_sc_hd__nor2_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18440_ _19619_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _15631_/A _15630_/B _15628_/X vssd1 vssd1 vccd1 vccd1 _15653_/B sky130_fd_sc_hd__a21o_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _13303_/B2 _12848_/X _12863_/X vssd1 vssd1 vccd1 vccd1 _13978_/B sky130_fd_sc_hd__a21oi_4
XFILLER_233_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14603_ _16595_/A0 _18410_/Q _14631_/S vssd1 vssd1 vccd1 vccd1 _18410_/D sky130_fd_sc_hd__mux2_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18371_ _19155_/CLK _18371_/D vssd1 vssd1 vccd1 vccd1 _18371_/Q sky130_fd_sc_hd__dfxtp_1
X_11815_ _11865_/A wire989/X vssd1 vssd1 vccd1 vccd1 _11815_/Y sky130_fd_sc_hd__nor2_4
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _15621_/C _15583_/B vssd1 vssd1 vccd1 vccd1 _15583_/Y sky130_fd_sc_hd__nor2_1
X_12795_ _12793_/X _12794_/X _12943_/S vssd1 vssd1 vccd1 vccd1 _12795_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17322_/A _17322_/B vssd1 vssd1 vccd1 vccd1 _19458_/D sky130_fd_sc_hd__and2_1
XFILLER_159_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14534_ _14596_/A _14534_/B vssd1 vssd1 vccd1 vccd1 _18375_/D sky130_fd_sc_hd__or2_1
X_11746_ _11746_/A _13127_/A vssd1 vssd1 vccd1 vccd1 _13125_/A sky130_fd_sc_hd__xnor2_4
XFILLER_144_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17253_ _17448_/A _17250_/B _18112_/Q _17389_/B1 vssd1 vssd1 vccd1 vccd1 _17253_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14465_ _18317_/Q _16470_/A0 _14485_/S vssd1 vssd1 vccd1 vccd1 _18317_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ _13465_/A _11677_/B vssd1 vssd1 vccd1 vccd1 _13476_/B sky130_fd_sc_hd__xnor2_4
XFILLER_128_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16204_ _16204_/A0 _18820_/Q _16222_/S vssd1 vssd1 vccd1 vccd1 _18820_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13416_ _13136_/S _12751_/Y _13414_/Y _13415_/Y vssd1 vssd1 vccd1 vccd1 _13416_/X
+ sky130_fd_sc_hd__a22o_2
X_10628_ _10633_/A _10627_/X _11563_/B1 vssd1 vssd1 vccd1 vccd1 _10628_/X sky130_fd_sc_hd__o21a_1
X_14396_ _16471_/A0 _18247_/Q _14415_/S vssd1 vssd1 vccd1 vccd1 _18247_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17184_ _17202_/A _17184_/B vssd1 vssd1 vccd1 vccd1 _17498_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16135_ _18770_/Q _16141_/B vssd1 vssd1 vccd1 vccd1 _16135_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13347_ _13438_/A _13333_/Y _13956_/B1 vssd1 vssd1 vccd1 vccd1 _13347_/X sky130_fd_sc_hd__a21o_1
X_10559_ _18650_/Q _18072_/Q _19091_/Q _18995_/Q _09108_/B _11559_/S1 vssd1 vssd1
+ vccd1 vccd1 _10559_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13278_ _19403_/Q _12579_/Y _12771_/X _13277_/X _12581_/Y vssd1 vssd1 vccd1 vccd1
+ _13278_/X sky130_fd_sc_hd__a221o_1
X_16066_ _18740_/Q _16054_/A _16069_/A _15845_/A vssd1 vssd1 vccd1 vccd1 _16066_/X
+ sky130_fd_sc_hd__a31o_1
X_12229_ _17875_/Q _12232_/C _12241_/A vssd1 vssd1 vccd1 vccd1 _12229_/Y sky130_fd_sc_hd__a21oi_1
X_15017_ _18506_/Q input206/X _16627_/S vssd1 vssd1 vccd1 vccd1 _18506_/D sky130_fd_sc_hd__mux2_1
XFILLER_64_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16968_ _16968_/A _16968_/B vssd1 vssd1 vccd1 vccd1 _19326_/D sky130_fd_sc_hd__and2_1
XFILLER_65_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18707_ _19306_/CLK _18707_/D vssd1 vssd1 vccd1 vccd1 _18707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15919_ _18682_/Q _15943_/A2 _15918_/X _15946_/C1 vssd1 vssd1 vccd1 vccd1 _18682_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16899_ _19309_/Q _17585_/A _16963_/S vssd1 vssd1 vccd1 vccd1 _16900_/B sky130_fd_sc_hd__mux2_1
XFILLER_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09440_ _18633_/Q _18055_/Q _09671_/S vssd1 vssd1 vccd1 vccd1 _09440_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18638_ _19142_/CLK _18638_/D vssd1 vssd1 vccd1 vccd1 _18638_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_65_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09371_ _10294_/A1 _18141_/Q _18787_/Q _09704_/S _10293_/B1 vssd1 vssd1 vccd1 vccd1
+ _09371_/X sky130_fd_sc_hd__a221o_1
XFILLER_52_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18569_ _19399_/CLK _18569_/D vssd1 vssd1 vccd1 vccd1 _18569_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_178_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput285 _11960_/X vssd1 vssd1 vccd1 vccd1 addr0[0] sky130_fd_sc_hd__buf_4
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput296 _11912_/X vssd1 vssd1 vccd1 vccd1 addr1[2] sky130_fd_sc_hd__buf_4
XFILLER_0_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09707_ _10297_/A1 _09700_/X _09701_/X vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__o21ai_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09638_ _09636_/X _09637_/X _11161_/S vssd1 vssd1 vccd1 vccd1 _09639_/B sky130_fd_sc_hd__mux2_1
XFILLER_216_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09569_ input128/X input164/X _09655_/S vssd1 vssd1 vccd1 vccd1 _09569_/X sky130_fd_sc_hd__mux2_8
XFILLER_215_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11600_ _10663_/S _11595_/X _11596_/X vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__o21ai_1
XFILLER_12_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ _12580_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _12580_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11531_ _13485_/A _11676_/B _13487_/S vssd1 vssd1 vccd1 vccd1 _11675_/B sky130_fd_sc_hd__a21oi_4
XFILLER_157_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14250_ _18123_/Q _14260_/B vssd1 vssd1 vccd1 vccd1 _14250_/X sky130_fd_sc_hd__or2_1
X_11462_ _18028_/Q _17996_/Q _11462_/S vssd1 vssd1 vccd1 vccd1 _11462_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13201_ _18110_/Q _13201_/B vssd1 vssd1 vccd1 vccd1 _13202_/B sky130_fd_sc_hd__nor2_1
XFILLER_171_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10413_ _10399_/A _10412_/Y _10399_/Y _11333_/A1 vssd1 vssd1 vccd1 vccd1 _10413_/Y
+ sky130_fd_sc_hd__o211ai_4
X_14181_ _14181_/A _14181_/B vssd1 vssd1 vccd1 vccd1 _18088_/D sky130_fd_sc_hd__and2_1
XFILLER_99_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11393_ _11391_/X _11392_/X _11478_/S vssd1 vssd1 vccd1 vccd1 _11393_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13132_ _13130_/A _12942_/X _13354_/A vssd1 vssd1 vccd1 vccd1 _13132_/X sky130_fd_sc_hd__a21o_1
X_10344_ _18334_/Q _17785_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _10344_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17940_ _18700_/CLK _17940_/D vssd1 vssd1 vccd1 vccd1 _17940_/Q sky130_fd_sc_hd__dfxtp_2
X_13063_ _19430_/Q _12560_/B _12560_/A vssd1 vssd1 vccd1 vccd1 _13063_/X sky130_fd_sc_hd__o21a_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10275_ _10273_/X _10274_/X _10275_/S vssd1 vssd1 vccd1 vccd1 _10275_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1400 fanout1407/X vssd1 vssd1 vccd1 vccd1 _09937_/S sky130_fd_sc_hd__buf_4
X_12014_ _17781_/Q _17682_/A0 _12022_/S vssd1 vssd1 vccd1 vccd1 _17781_/D sky130_fd_sc_hd__mux2_1
Xfanout1411 fanout1415/X vssd1 vssd1 vccd1 vccd1 _09344_/S sky130_fd_sc_hd__buf_4
XFILLER_151_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1422 _11403_/S vssd1 vssd1 vccd1 vccd1 _11384_/B sky130_fd_sc_hd__buf_2
X_17871_ _19310_/CLK _17871_/D vssd1 vssd1 vccd1 vccd1 _17871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1433 _10009_/A vssd1 vssd1 vccd1 vccd1 _11484_/B1 sky130_fd_sc_hd__buf_12
Xfanout1444 _10408_/S vssd1 vssd1 vccd1 vccd1 _10403_/S sky130_fd_sc_hd__buf_6
X_19610_ _19638_/CLK _19610_/D vssd1 vssd1 vccd1 vccd1 _19610_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1455 _09136_/S vssd1 vssd1 vccd1 vccd1 _11464_/C1 sky130_fd_sc_hd__buf_6
X_16822_ _16839_/A _16839_/B _16840_/B vssd1 vssd1 vccd1 vccd1 _16824_/A sky130_fd_sc_hd__and3_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1466 fanout1469/X vssd1 vssd1 vccd1 vccd1 _11353_/B2 sky130_fd_sc_hd__buf_4
XFILLER_66_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1477 _09801_/S vssd1 vssd1 vccd1 vccd1 _11125_/B2 sky130_fd_sc_hd__buf_6
XFILLER_254_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout490 _14889_/B1 vssd1 vssd1 vccd1 vccd1 _15010_/B1 sky130_fd_sc_hd__buf_12
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1488 _10496_/B vssd1 vssd1 vccd1 vccd1 _09885_/S sky130_fd_sc_hd__buf_4
XFILLER_219_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1499 fanout1525/X vssd1 vssd1 vccd1 vccd1 _10290_/S sky130_fd_sc_hd__buf_4
X_19541_ _19553_/CLK _19541_/D vssd1 vssd1 vccd1 vccd1 _19541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16753_ _19271_/Q _16754_/B vssd1 vssd1 vccd1 vccd1 _16755_/B sky130_fd_sc_hd__nor2_1
XFILLER_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13965_ _12656_/B _12837_/B _14154_/B1 _12739_/X _13964_/Y vssd1 vssd1 vccd1 vccd1
+ _13965_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15704_ _18589_/Q _18588_/Q _15704_/C vssd1 vssd1 vccd1 vccd1 _15746_/C sky130_fd_sc_hd__and3_2
XFILLER_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12916_ _19299_/Q _12583_/Y _12914_/X _12915_/X vssd1 vssd1 vccd1 vccd1 _12916_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19472_ _19543_/CLK _19472_/D vssd1 vssd1 vccd1 vccd1 _19472_/Q sky130_fd_sc_hd__dfxtp_1
X_16684_ _19247_/Q _16675_/C _16678_/Y vssd1 vssd1 vccd1 vccd1 _19247_/D sky130_fd_sc_hd__o21a_1
XFILLER_250_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13896_ _12712_/S _12891_/X _12897_/X _13896_/B2 vssd1 vssd1 vccd1 vccd1 _13896_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_261_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18423_ _19197_/CLK _18423_/D vssd1 vssd1 vccd1 vccd1 _18423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15635_ _13737_/X _15110_/X _10599_/Y _15111_/A vssd1 vssd1 vccd1 vccd1 _15635_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _15481_/A _15130_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _12847_/X sky130_fd_sc_hd__mux2_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18354_ _19632_/CLK _18354_/D vssd1 vssd1 vccd1 vccd1 _18354_/Q sky130_fd_sc_hd__dfxtp_1
X_15566_ _19476_/Q _19410_/Q vssd1 vssd1 vccd1 vccd1 _15568_/A sky130_fd_sc_hd__nand2_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12770_/X _12777_/X _12859_/S vssd1 vssd1 vccd1 vccd1 _12778_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _18129_/Q _15782_/A1 _17205_/Y _17307_/B vssd1 vssd1 vccd1 vccd1 _17305_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14517_ _16619_/A0 _18367_/Q _14517_/S vssd1 vssd1 vccd1 vccd1 _18367_/D sky130_fd_sc_hd__mux2_1
X_18285_ _18741_/CLK _18285_/D vssd1 vssd1 vccd1 vccd1 _18285_/Q sky130_fd_sc_hd__dfxtp_1
X_11729_ _11726_/B _15039_/B vssd1 vssd1 vccd1 vccd1 _11729_/X sky130_fd_sc_hd__and2b_2
X_15497_ _15497_/A _15497_/B vssd1 vssd1 vccd1 vccd1 _15497_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_175_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17236_ _18106_/Q _17382_/A _17418_/A _17256_/B vssd1 vssd1 vccd1 vccd1 _17236_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14448_ _18587_/Q _14450_/B vssd1 vssd1 vccd1 vccd1 _18300_/D sky130_fd_sc_hd__and2_1
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17167_ _19407_/Q fanout534/X _17468_/A _17212_/B2 vssd1 vssd1 vccd1 vccd1 _17168_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14379_ _18231_/Q _16553_/A0 _14382_/S vssd1 vssd1 vccd1 vccd1 _18231_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16118_ _16140_/A1 _16117_/Y _12107_/A vssd1 vssd1 vccd1 vccd1 _18761_/D sky130_fd_sc_hd__a21oi_1
XFILLER_155_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ _17187_/B _17116_/A2 _17097_/X _17592_/B vssd1 vssd1 vccd1 vccd1 _19382_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08940_ _12029_/A _08940_/B vssd1 vssd1 vccd1 vccd1 _08940_/X sky130_fd_sc_hd__or2_4
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16049_ _18729_/Q _18736_/Q _16051_/S vssd1 vssd1 vccd1 vccd1 _16050_/B sky130_fd_sc_hd__mux2_1
XFILLER_131_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08871_ _17898_/Q _17897_/Q _17896_/Q _17895_/Q vssd1 vssd1 vccd1 vccd1 _08872_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09423_ _10300_/S _09422_/X _11495_/B1 vssd1 vssd1 vccd1 vccd1 _09424_/B sky130_fd_sc_hd__a21o_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09354_ _18056_/Q _10101_/B _09353_/X _10335_/S vssd1 vssd1 vccd1 vccd1 _09354_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09285_ _09494_/A _18820_/Q _09285_/C vssd1 vssd1 vccd1 vccd1 _09285_/X sky130_fd_sc_hd__and3_1
XFILLER_138_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_148_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19525_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ _10043_/X _10044_/Y _10059_/X _11279_/B1 vssd1 vssd1 vccd1 vccd1 _10060_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13750_ _19417_/Q _13948_/A2 _13948_/B1 vssd1 vssd1 vccd1 vccd1 _13750_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10962_ _10040_/S _10961_/X _11623_/A1 vssd1 vssd1 vccd1 vccd1 _10963_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ _12685_/X _12700_/X _13135_/S vssd1 vssd1 vccd1 vccd1 _12702_/A sky130_fd_sc_hd__mux2_2
X_13681_ _19255_/Q _13943_/A2 _13943_/B1 _19287_/Q vssd1 vssd1 vccd1 vccd1 _13681_/X
+ sky130_fd_sc_hd__a22o_2
X_10893_ _11606_/S _10890_/X _10892_/X vssd1 vssd1 vccd1 vccd1 _10901_/B sky130_fd_sc_hd__a21oi_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15420_ _15399_/A _15398_/B _15398_/A vssd1 vssd1 vccd1 vccd1 _15421_/B sky130_fd_sc_hd__a21boi_2
XPHY_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12632_ _13485_/A _11214_/A _11212_/Y _11136_/Y _11138_/A vssd1 vssd1 vccd1 vccd1
+ _12632_/X sky130_fd_sc_hd__o32a_1
XPHY_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12563_ _12563_/A _12563_/B vssd1 vssd1 vccd1 vccd1 _13167_/B sky130_fd_sc_hd__or2_4
X_15351_ _18573_/Q _15351_/A2 _15350_/Y _17469_/C1 vssd1 vssd1 vccd1 vccd1 _18573_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_200_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11514_ _11512_/X _11513_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _11514_/X sky130_fd_sc_hd__mux2_1
X_14302_ _16455_/A1 _18161_/Q _14304_/S vssd1 vssd1 vccd1 vccd1 _18161_/D sky130_fd_sc_hd__mux2_1
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18070_ _19211_/CLK _18070_/D vssd1 vssd1 vccd1 vccd1 _18070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12494_ _12548_/A _12554_/B vssd1 vssd1 vccd1 vccd1 _12544_/A sky130_fd_sc_hd__or2_4
XFILLER_157_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15282_ _17389_/B1 _15281_/X _15274_/X _15424_/C1 vssd1 vssd1 vccd1 vccd1 _15282_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17021_ _19347_/Q _17041_/B vssd1 vssd1 vccd1 vccd1 _17021_/X sky130_fd_sc_hd__or2_1
X_14233_ _18288_/Q _14261_/A2 _14232_/X _14450_/B vssd1 vssd1 vccd1 vccd1 _18114_/D
+ sky130_fd_sc_hd__o211a_1
X_11445_ _12597_/A _11445_/B vssd1 vssd1 vccd1 vccd1 _11446_/B sky130_fd_sc_hd__nor2_4
XFILLER_153_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ _18720_/Q _14164_/B _15953_/A vssd1 vssd1 vccd1 vccd1 _16145_/B sky130_fd_sc_hd__or3_1
XFILLER_171_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11376_ _11452_/A _11376_/B vssd1 vssd1 vccd1 vccd1 _11376_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10327_ _18559_/Q _18434_/Q _18043_/Q _18011_/Q _09181_/S _11001_/C1 vssd1 vssd1
+ vccd1 vccd1 _10327_/X sky130_fd_sc_hd__mux4_1
X_13115_ _17862_/Q _13945_/A2 _13104_/X _13115_/B2 _13115_/C1 vssd1 vssd1 vccd1 vccd1
+ _13116_/B sky130_fd_sc_hd__a221o_1
X_18972_ _19624_/CLK _18972_/D vssd1 vssd1 vccd1 vccd1 _18972_/Q sky130_fd_sc_hd__dfxtp_1
X_14095_ _17678_/A0 _18035_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _18035_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17923_ _18201_/CLK _17923_/D vssd1 vssd1 vccd1 vccd1 _17923_/Q sky130_fd_sc_hd__dfxtp_4
X_13046_ _13046_/A1 _12883_/A _12745_/X vssd1 vssd1 vccd1 vccd1 _13047_/A sky130_fd_sc_hd__o21a_1
X_10258_ _10263_/A1 _17786_/Q _10253_/C _18335_/Q vssd1 vssd1 vccd1 vccd1 _10258_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1230 _14692_/A2 vssd1 vssd1 vccd1 vccd1 _14934_/C sky130_fd_sc_hd__buf_6
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1241 _09108_/X vssd1 vssd1 vccd1 vccd1 _11023_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_267_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17854_ _19268_/CLK _17854_/D vssd1 vssd1 vccd1 vccd1 _17854_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ _10187_/X _10188_/X _10335_/S vssd1 vssd1 vccd1 vccd1 _10190_/B sky130_fd_sc_hd__mux2_1
Xfanout1252 _11337_/B vssd1 vssd1 vccd1 vccd1 _11135_/S sky130_fd_sc_hd__buf_6
XFILLER_282_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1263 _08890_/Y vssd1 vssd1 vccd1 vccd1 _09141_/A sky130_fd_sc_hd__buf_12
XFILLER_227_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1274 _12264_/X vssd1 vssd1 vccd1 vccd1 _14153_/A sky130_fd_sc_hd__buf_6
Xfanout1285 _15970_/A2 vssd1 vssd1 vccd1 vccd1 _16002_/A2 sky130_fd_sc_hd__buf_4
X_16805_ _19290_/Q _16807_/C _16804_/Y vssd1 vssd1 vccd1 vccd1 _19290_/D sky130_fd_sc_hd__a21oi_1
XFILLER_282_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1296 _14586_/A vssd1 vssd1 vccd1 vccd1 _14592_/A sky130_fd_sc_hd__clkbuf_4
X_17785_ _19613_/CLK _17785_/D vssd1 vssd1 vccd1 vccd1 _17785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14997_ input66/X input101/X _15007_/S vssd1 vssd1 vccd1 vccd1 _14998_/A sky130_fd_sc_hd__mux2_2
XFILLER_47_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19524_ _19526_/CLK _19524_/D vssd1 vssd1 vccd1 vccd1 _19524_/Q sky130_fd_sc_hd__dfxtp_1
X_16736_ _19265_/Q _19264_/Q _19263_/Q _16736_/D vssd1 vssd1 vccd1 vccd1 _16743_/C
+ sky130_fd_sc_hd__and4_1
X_13948_ _19423_/Q _13948_/A2 _13948_/B1 vssd1 vssd1 vccd1 vccd1 _13948_/X sky130_fd_sc_hd__a21o_1
XFILLER_90_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19455_ _19521_/CLK _19455_/D vssd1 vssd1 vccd1 vccd1 _19455_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16667_ _19244_/Q _19243_/Q _16667_/C vssd1 vssd1 vccd1 vccd1 _16674_/C sky130_fd_sc_hd__and3_1
XFILLER_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13879_ _19551_/Q _13946_/B vssd1 vssd1 vccd1 vccd1 _13879_/X sky130_fd_sc_hd__or2_1
XFILLER_250_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18406_ _19477_/CLK _18406_/D vssd1 vssd1 vccd1 vccd1 _18406_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_201_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15618_ _15702_/A _15618_/B vssd1 vssd1 vccd1 vccd1 _15638_/D sky130_fd_sc_hd__xnor2_1
X_19386_ _19481_/CLK _19386_/D vssd1 vssd1 vccd1 vccd1 _19386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16598_ _17665_/A0 _19201_/Q _16619_/S vssd1 vssd1 vccd1 vccd1 _19201_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18337_ _19615_/CLK _18337_/D vssd1 vssd1 vccd1 vccd1 _18337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15549_ _15549_/A _15623_/A vssd1 vssd1 vccd1 vccd1 _15702_/A sky130_fd_sc_hd__nand2_8
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09070_ _17894_/Q _17893_/Q _12443_/A _09070_/D vssd1 vssd1 vccd1 vccd1 _12740_/A
+ sky130_fd_sc_hd__or4_2
X_18268_ _18973_/CLK _18268_/D vssd1 vssd1 vccd1 vccd1 _18268_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17219_ _17219_/A _17219_/B vssd1 vssd1 vccd1 vccd1 _17219_/Y sky130_fd_sc_hd__nor2_2
XFILLER_162_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18199_ _18201_/CLK _18199_/D vssd1 vssd1 vccd1 vccd1 _18199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09972_ _09970_/X _09971_/X _09972_/S vssd1 vssd1 vccd1 vccd1 _09972_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08923_ _12089_/A _17798_/Q vssd1 vssd1 vccd1 vccd1 _14074_/B sky130_fd_sc_hd__nand2_4
XFILLER_131_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08854_ _17894_/Q vssd1 vssd1 vccd1 vccd1 _08870_/A sky130_fd_sc_hd__inv_2
XFILLER_285_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09406_ _18539_/Q _18414_/Q _18023_/Q _17991_/Q _09428_/B2 _11199_/S1 vssd1 vssd1
+ vccd1 vccd1 _09406_/X sky130_fd_sc_hd__mux4_1
XFILLER_240_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09337_ _09335_/X _09336_/X _10265_/A vssd1 vssd1 vccd1 vccd1 _09337_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09268_ _18057_/Q _11479_/B _09267_/X _10408_/S vssd1 vssd1 vccd1 vccd1 _09268_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ _18853_/Q _18885_/Q _10141_/S vssd1 vssd1 vccd1 vccd1 _09199_/X sky130_fd_sc_hd__mux2_1
XFILLER_267_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ _11568_/A _11228_/X _11229_/X _09099_/Y vssd1 vssd1 vccd1 vccd1 _11230_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11161_ _11159_/X _11160_/X _11161_/S vssd1 vssd1 vccd1 vccd1 _11161_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10112_ _11017_/A1 _18234_/Q _10176_/S _18969_/Q vssd1 vssd1 vccd1 vccd1 _10112_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_161_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ _11305_/A1 _18611_/Q _18182_/Q _11309_/S vssd1 vssd1 vccd1 vccd1 _11092_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14920_ _18493_/Q _15011_/A2 _14919_/Y _16787_/A vssd1 vssd1 vccd1 vccd1 _18493_/D
+ sky130_fd_sc_hd__a211o_1
X_10043_ _10589_/S _10042_/Y _10041_/Y _15481_/A vssd1 vssd1 vccd1 vccd1 _10043_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ _14849_/X _14850_/X _14714_/B vssd1 vssd1 vccd1 vccd1 _14851_/X sky130_fd_sc_hd__a21o_1
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _18127_/Q _18126_/Q _13802_/C vssd1 vssd1 vccd1 vccd1 _13837_/B sky130_fd_sc_hd__and3_1
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _19527_/Q _17561_/B _17588_/B1 _17569_/X vssd1 vssd1 vccd1 vccd1 _19527_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14782_ _18110_/Q _14994_/B _14771_/X _14781_/X vssd1 vssd1 vccd1 vccd1 _14782_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11994_ _17761_/Q _16595_/A0 _12022_/S vssd1 vssd1 vccd1 vccd1 _17761_/D sky130_fd_sc_hd__mux2_1
XFILLER_216_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16521_ _10239_/B _19127_/Q _16521_/S vssd1 vssd1 vccd1 vccd1 _19127_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13733_ _13966_/C1 _13731_/X _13732_/X _13729_/X vssd1 vssd1 vccd1 vccd1 _13733_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_232_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10945_ _10924_/X _10927_/X _10944_/X vssd1 vssd1 vccd1 vccd1 _10945_/X sky130_fd_sc_hd__a21o_1
XFILLER_188_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19653_/A
+ sky130_fd_sc_hd__clkbuf_16
X_19240_ _19273_/CLK _19240_/D vssd1 vssd1 vccd1 vccd1 _19240_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_188_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16452_ _19060_/Q _16617_/A0 _16453_/S vssd1 vssd1 vccd1 vccd1 _19060_/D sky130_fd_sc_hd__mux2_1
X_13664_ _13616_/A _13615_/A _12643_/B vssd1 vssd1 vccd1 vccd1 _13665_/B sky130_fd_sc_hd__o21ba_2
X_10876_ _11112_/A _10876_/B vssd1 vssd1 vccd1 vccd1 _10876_/Y sky130_fd_sc_hd__nand2_1
XFILLER_204_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15403_ _12755_/A _15429_/A2 _15484_/A vssd1 vssd1 vccd1 vccd1 _15408_/A sky130_fd_sc_hd__o21ai_4
X_19171_ _19203_/CLK _19171_/D vssd1 vssd1 vccd1 vccd1 _19171_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _12615_/A _12985_/B _12985_/A _13033_/A vssd1 vssd1 vccd1 vccd1 _13148_/B
+ sky130_fd_sc_hd__or4bb_2
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16383_ _16549_/A0 _18994_/Q _16391_/S vssd1 vssd1 vccd1 vccd1 _18994_/D sky130_fd_sc_hd__mux2_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _13637_/A _14014_/B _13581_/X vssd1 vssd1 vccd1 vccd1 _13595_/Y sky130_fd_sc_hd__o21ai_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18122_ _19453_/CLK _18122_/D vssd1 vssd1 vccd1 vccd1 _18122_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15334_ _18112_/Q _15133_/Y _15333_/X _15382_/B2 vssd1 vssd1 vccd1 vccd1 _15335_/B
+ sky130_fd_sc_hd__a22oi_2
X_12546_ _19232_/Q _13625_/A2 _13625_/B1 _19264_/Q vssd1 vssd1 vccd1 vccd1 _12546_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18053_ _19622_/CLK _18053_/D vssd1 vssd1 vccd1 vccd1 _18053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15265_ _15198_/X _15201_/X _15263_/C _15263_/D _15264_/Y vssd1 vssd1 vccd1 vccd1
+ _15265_/X sky130_fd_sc_hd__a41o_1
X_12477_ _12488_/A _17917_/Q _12476_/Y vssd1 vssd1 vccd1 vccd1 _12501_/B sky130_fd_sc_hd__a21o_1
XANTENNA_4 _18199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ _17579_/A _17008_/A2 _17003_/X _17338_/A vssd1 vssd1 vccd1 vccd1 _19338_/D
+ sky130_fd_sc_hd__o211a_1
X_14216_ _18106_/Q _14244_/B vssd1 vssd1 vccd1 vccd1 _14216_/X sky130_fd_sc_hd__or2_1
X_11428_ _11428_/A _11428_/B vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__and2_1
XFILLER_172_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15196_ _18106_/Q _15133_/Y _15195_/X _15216_/A1 vssd1 vssd1 vccd1 vccd1 _15199_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ _11360_/A1 _19632_/Q _18921_/Q _11360_/B2 vssd1 vssd1 vccd1 vccd1 _11359_/X
+ sky130_fd_sc_hd__a22o_1
X_14147_ _14147_/A _14147_/B _14147_/C _14147_/D vssd1 vssd1 vccd1 vccd1 _14149_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18955_ _19147_/CLK _18955_/D vssd1 vssd1 vccd1 vccd1 _18955_/Q sky130_fd_sc_hd__dfxtp_1
X_14078_ _17694_/A0 _18018_/Q _14098_/S vssd1 vssd1 vccd1 vccd1 _18018_/D sky130_fd_sc_hd__mux2_1
XFILLER_258_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17906_ _18817_/CLK _17906_/D vssd1 vssd1 vccd1 vccd1 _17906_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13029_ _14214_/A _13028_/C _18106_/Q vssd1 vssd1 vccd1 vccd1 _13030_/B sky130_fd_sc_hd__a21oi_1
XFILLER_255_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18886_ _19206_/CLK _18886_/D vssd1 vssd1 vccd1 vccd1 _18886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1060 _13483_/B vssd1 vssd1 vccd1 vccd1 _13961_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_266_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1071 _14027_/A2 vssd1 vssd1 vccd1 vccd1 _14004_/A sky130_fd_sc_hd__buf_6
XFILLER_255_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17837_ _19310_/CLK _17837_/D vssd1 vssd1 vccd1 vccd1 _17837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1082 _09980_/A2 vssd1 vssd1 vccd1 vccd1 _16593_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_187_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1093 _09697_/B vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__buf_6
XFILLER_254_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17768_ _19596_/CLK _17768_/D vssd1 vssd1 vccd1 vccd1 _17768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16719_ _19259_/Q _16723_/C _16964_/A vssd1 vssd1 vccd1 vccd1 _16719_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_223_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19507_ _19507_/CLK _19507_/D vssd1 vssd1 vccd1 vccd1 _19507_/Q sky130_fd_sc_hd__dfxtp_1
X_17699_ _17699_/A0 _19625_/Q _17719_/S vssd1 vssd1 vccd1 vccd1 _19625_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19438_ _19552_/CLK _19438_/D vssd1 vssd1 vccd1 vccd1 _19438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19369_ _19465_/CLK _19369_/D vssd1 vssd1 vccd1 vccd1 _19369_/Q sky130_fd_sc_hd__dfxtp_1
X_09122_ _11465_/A1 _19565_/Q _11455_/S _19597_/Q _09135_/S vssd1 vssd1 vccd1 vccd1
+ _09122_/X sky130_fd_sc_hd__o221a_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _17963_/Q _11295_/A2 _08947_/A _17931_/Q _08946_/B vssd1 vssd1 vccd1 vccd1
+ _09053_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_191_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09955_ _18844_/Q _09952_/S _10144_/B1 vssd1 vssd1 vccd1 vccd1 _09955_/X sky130_fd_sc_hd__o21a_1
XFILLER_103_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08906_ _08932_/A _12053_/A _17802_/Q _12051_/A vssd1 vssd1 vccd1 vccd1 _11556_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_103_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09886_ _10033_/S _09885_/X _09884_/X _11274_/S1 vssd1 vssd1 vccd1 vccd1 _09886_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08837_ _09245_/A vssd1 vssd1 vccd1 vccd1 _08837_/Y sky130_fd_sc_hd__clkinv_2
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_405 _13818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_416 _13647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_427 _11822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_438 _13986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_449 _13757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10730_ _11622_/A1 _10719_/X _10729_/X _08950_/A vssd1 vssd1 vccd1 vccd1 _10730_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10661_ _18866_/Q _18898_/Q _10667_/S vssd1 vssd1 vccd1 vccd1 _10661_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ _12412_/A _12400_/B vssd1 vssd1 vccd1 vccd1 _12400_/Y sky130_fd_sc_hd__nand2_1
X_13380_ _17837_/Q _13821_/B _13379_/X vssd1 vssd1 vccd1 vccd1 _13380_/X sky130_fd_sc_hd__o21a_1
XFILLER_185_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10592_ _19642_/Q _18931_/Q _10667_/S vssd1 vssd1 vccd1 vccd1 _10592_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _17807_/Q _17806_/Q _17805_/Q _17804_/Q vssd1 vssd1 vccd1 vccd1 _12332_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_182_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_163_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19553_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12262_ _12443_/A _12315_/B _12665_/B vssd1 vssd1 vccd1 vccd1 _12263_/A sky130_fd_sc_hd__or3b_4
X_15050_ _18534_/Q _17694_/A0 _15070_/S vssd1 vssd1 vccd1 vccd1 _18534_/D sky130_fd_sc_hd__mux2_1
X_14001_ _17965_/Q _14034_/B _14000_/Y _14001_/C1 vssd1 vssd1 vccd1 vccd1 _17965_/D
+ sky130_fd_sc_hd__o211a_1
X_11213_ _11214_/A _11214_/B vssd1 vssd1 vccd1 vccd1 _13468_/S sky130_fd_sc_hd__and2_2
XFILLER_269_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12193_ _16752_/A _12193_/B _12194_/B vssd1 vssd1 vccd1 vccd1 _17861_/D sky130_fd_sc_hd__nor3_1
XFILLER_150_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11144_ _17936_/Q _08948_/B _11143_/X _08947_/B vssd1 vssd1 vccd1 vccd1 _11144_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18740_ _18741_/CLK _18740_/D vssd1 vssd1 vccd1 vccd1 _18740_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15952_ _15951_/X _15952_/B vssd1 vssd1 vccd1 vccd1 _18693_/D sky130_fd_sc_hd__and2b_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11075_ _18549_/Q _11094_/S vssd1 vssd1 vccd1 vccd1 _11075_/X sky130_fd_sc_hd__or2_1
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput130 dout1[30] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_hd__clkbuf_2
XFILLER_283_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput141 dout1[40] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_hd__buf_2
Xinput152 dout1[50] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_hd__buf_2
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10026_ _15120_/A _11782_/B _10025_/Y _10027_/B vssd1 vssd1 vccd1 vccd1 _10026_/X
+ sky130_fd_sc_hd__a211o_1
X_14903_ _14901_/X _14902_/X _14714_/B vssd1 vssd1 vccd1 vccd1 _14903_/X sky130_fd_sc_hd__a21o_1
Xinput163 dout1[60] vssd1 vssd1 vccd1 vccd1 input163/X sky130_fd_sc_hd__buf_2
X_18671_ _18683_/CLK _18671_/D vssd1 vssd1 vccd1 vccd1 _18671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15883_ _18670_/Q _15949_/A2 _15882_/X _15904_/C1 vssd1 vssd1 vccd1 vccd1 _18670_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput174 irq[12] vssd1 vssd1 vccd1 vccd1 _15089_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_37_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput185 irq[8] vssd1 vssd1 vccd1 vccd1 input185/X sky130_fd_sc_hd__buf_2
XFILLER_252_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput196 localMemory_wb_adr_i[15] vssd1 vssd1 vccd1 vccd1 input196/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17622_ _19552_/Q _17622_/A2 _17621_/X _17352_/A vssd1 vssd1 vccd1 vccd1 _19552_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ input48/X input83/X _14844_/S vssd1 vssd1 vccd1 vccd1 _14835_/A sky130_fd_sc_hd__mux2_1
XFILLER_264_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _17214_/Y _17493_/B _17552_/X _16048_/A vssd1 vssd1 vccd1 vccd1 _17553_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_251_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _14718_/A _14764_/X _14846_/B1 vssd1 vssd1 vccd1 vccd1 _14765_/Y sky130_fd_sc_hd__o21bai_4
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ _15845_/B _11977_/B _18692_/Q vssd1 vssd1 vccd1 vccd1 _11977_/X sky130_fd_sc_hd__or3b_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16504_ _17670_/A0 _19110_/Q _16523_/S vssd1 vssd1 vccd1 vccd1 _19110_/D sky130_fd_sc_hd__mux2_1
X_13716_ _19546_/Q _13921_/S vssd1 vssd1 vccd1 vccd1 _13716_/X sky130_fd_sc_hd__or2_1
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10928_ _18458_/Q _18359_/Q _10940_/S vssd1 vssd1 vccd1 vccd1 _10928_/X sky130_fd_sc_hd__mux2_1
X_17484_ _19508_/Q _17523_/B _17482_/X _17483_/Y _17354_/A vssd1 vssd1 vccd1 vccd1
+ _19508_/D sky130_fd_sc_hd__o221a_1
XFILLER_220_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14696_ _14696_/A _18269_/Q vssd1 vssd1 vccd1 vccd1 _14718_/A sky130_fd_sc_hd__nand2_8
XFILLER_32_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19223_ _19625_/CLK _19223_/D vssd1 vssd1 vccd1 vccd1 _19223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16435_ _19043_/Q _17667_/A0 _16457_/S vssd1 vssd1 vccd1 vccd1 _19043_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13647_ _13647_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13647_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10859_ _11328_/S _10854_/X _10858_/X _11579_/A vssd1 vssd1 vccd1 vccd1 _10859_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_258_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19154_ _19154_/CLK _19154_/D vssd1 vssd1 vccd1 vccd1 _19154_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16532_/A0 _18977_/Q _16385_/S vssd1 vssd1 vccd1 vccd1 _18977_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13938_/A _13566_/A _13971_/A2 _12320_/B vssd1 vssd1 vccd1 vccd1 _13579_/B
+ sky130_fd_sc_hd__a22o_1
X_18105_ _18734_/CLK _18105_/D vssd1 vssd1 vccd1 vccd1 _18105_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15317_ _19434_/Q _15411_/B _17211_/A _15316_/Y vssd1 vssd1 vccd1 vccd1 _15317_/Y
+ sky130_fd_sc_hd__o211ai_1
X_19085_ _19604_/CLK _19085_/D vssd1 vssd1 vccd1 vccd1 _19085_/Q sky130_fd_sc_hd__dfxtp_1
X_12529_ _12768_/A _13165_/C vssd1 vssd1 vccd1 vccd1 _12529_/Y sky130_fd_sc_hd__nor2_8
X_16297_ _17695_/A0 _18910_/Q _16320_/S vssd1 vssd1 vccd1 vccd1 _18910_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18036_ _19575_/CLK _18036_/D vssd1 vssd1 vccd1 vccd1 _18036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15248_ _15263_/D _15248_/B vssd1 vssd1 vccd1 vccd1 _15248_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_173_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _15179_/A _15179_/B vssd1 vssd1 vccd1 vccd1 _15179_/X sky130_fd_sc_hd__and2_1
XFILLER_125_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _11556_/C _09739_/X _11687_/A vssd1 vssd1 vccd1 vccd1 _09740_/X sky130_fd_sc_hd__o21a_1
X_18938_ _19649_/CLK _18938_/D vssd1 vssd1 vccd1 vccd1 _18938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
.ends

