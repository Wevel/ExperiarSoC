magic
tech sky130A
magscale 1 2
timestamp 1651534092
<< obsli1 >>
rect 1104 2159 108836 147441
<< obsm1 >>
rect 474 2128 109558 147552
<< metal2 >>
rect 478 149200 534 150000
rect 1398 149200 1454 150000
rect 2318 149200 2374 150000
rect 3330 149200 3386 150000
rect 4250 149200 4306 150000
rect 5262 149200 5318 150000
rect 6182 149200 6238 150000
rect 7194 149200 7250 150000
rect 8114 149200 8170 150000
rect 9126 149200 9182 150000
rect 10046 149200 10102 150000
rect 11058 149200 11114 150000
rect 11978 149200 12034 150000
rect 12990 149200 13046 150000
rect 13910 149200 13966 150000
rect 14922 149200 14978 150000
rect 15842 149200 15898 150000
rect 16854 149200 16910 150000
rect 17774 149200 17830 150000
rect 18786 149200 18842 150000
rect 19706 149200 19762 150000
rect 20718 149200 20774 150000
rect 21638 149200 21694 150000
rect 22650 149200 22706 150000
rect 23570 149200 23626 150000
rect 24582 149200 24638 150000
rect 25502 149200 25558 150000
rect 26514 149200 26570 150000
rect 27434 149200 27490 150000
rect 28446 149200 28502 150000
rect 29366 149200 29422 150000
rect 30378 149200 30434 150000
rect 31298 149200 31354 150000
rect 32310 149200 32366 150000
rect 33230 149200 33286 150000
rect 34242 149200 34298 150000
rect 35162 149200 35218 150000
rect 36174 149200 36230 150000
rect 37094 149200 37150 150000
rect 38106 149200 38162 150000
rect 39026 149200 39082 150000
rect 40038 149200 40094 150000
rect 40958 149200 41014 150000
rect 41970 149200 42026 150000
rect 42890 149200 42946 150000
rect 43902 149200 43958 150000
rect 44822 149200 44878 150000
rect 45834 149200 45890 150000
rect 46754 149200 46810 150000
rect 47766 149200 47822 150000
rect 48686 149200 48742 150000
rect 49698 149200 49754 150000
rect 50618 149200 50674 150000
rect 51630 149200 51686 150000
rect 52550 149200 52606 150000
rect 53562 149200 53618 150000
rect 54482 149200 54538 150000
rect 55494 149200 55550 150000
rect 56414 149200 56470 150000
rect 57334 149200 57390 150000
rect 58346 149200 58402 150000
rect 59266 149200 59322 150000
rect 60278 149200 60334 150000
rect 61198 149200 61254 150000
rect 62210 149200 62266 150000
rect 63130 149200 63186 150000
rect 64142 149200 64198 150000
rect 65062 149200 65118 150000
rect 66074 149200 66130 150000
rect 66994 149200 67050 150000
rect 68006 149200 68062 150000
rect 68926 149200 68982 150000
rect 69938 149200 69994 150000
rect 70858 149200 70914 150000
rect 71870 149200 71926 150000
rect 72790 149200 72846 150000
rect 73802 149200 73858 150000
rect 74722 149200 74778 150000
rect 75734 149200 75790 150000
rect 76654 149200 76710 150000
rect 77666 149200 77722 150000
rect 78586 149200 78642 150000
rect 79598 149200 79654 150000
rect 80518 149200 80574 150000
rect 81530 149200 81586 150000
rect 82450 149200 82506 150000
rect 83462 149200 83518 150000
rect 84382 149200 84438 150000
rect 85394 149200 85450 150000
rect 86314 149200 86370 150000
rect 87326 149200 87382 150000
rect 88246 149200 88302 150000
rect 89258 149200 89314 150000
rect 90178 149200 90234 150000
rect 91190 149200 91246 150000
rect 92110 149200 92166 150000
rect 93122 149200 93178 150000
rect 94042 149200 94098 150000
rect 95054 149200 95110 150000
rect 95974 149200 96030 150000
rect 96986 149200 97042 150000
rect 97906 149200 97962 150000
rect 98918 149200 98974 150000
rect 99838 149200 99894 150000
rect 100850 149200 100906 150000
rect 101770 149200 101826 150000
rect 102782 149200 102838 150000
rect 103702 149200 103758 150000
rect 104714 149200 104770 150000
rect 105634 149200 105690 150000
rect 106646 149200 106702 150000
rect 107566 149200 107622 150000
rect 108578 149200 108634 150000
rect 109498 149200 109554 150000
<< obsm2 >>
rect 590 149144 1342 149274
rect 1510 149144 2262 149274
rect 2430 149144 3274 149274
rect 3442 149144 4194 149274
rect 4362 149144 5206 149274
rect 5374 149144 6126 149274
rect 6294 149144 7138 149274
rect 7306 149144 8058 149274
rect 8226 149144 9070 149274
rect 9238 149144 9990 149274
rect 10158 149144 11002 149274
rect 11170 149144 11922 149274
rect 12090 149144 12934 149274
rect 13102 149144 13854 149274
rect 14022 149144 14866 149274
rect 15034 149144 15786 149274
rect 15954 149144 16798 149274
rect 16966 149144 17718 149274
rect 17886 149144 18730 149274
rect 18898 149144 19650 149274
rect 19818 149144 20662 149274
rect 20830 149144 21582 149274
rect 21750 149144 22594 149274
rect 22762 149144 23514 149274
rect 23682 149144 24526 149274
rect 24694 149144 25446 149274
rect 25614 149144 26458 149274
rect 26626 149144 27378 149274
rect 27546 149144 28390 149274
rect 28558 149144 29310 149274
rect 29478 149144 30322 149274
rect 30490 149144 31242 149274
rect 31410 149144 32254 149274
rect 32422 149144 33174 149274
rect 33342 149144 34186 149274
rect 34354 149144 35106 149274
rect 35274 149144 36118 149274
rect 36286 149144 37038 149274
rect 37206 149144 38050 149274
rect 38218 149144 38970 149274
rect 39138 149144 39982 149274
rect 40150 149144 40902 149274
rect 41070 149144 41914 149274
rect 42082 149144 42834 149274
rect 43002 149144 43846 149274
rect 44014 149144 44766 149274
rect 44934 149144 45778 149274
rect 45946 149144 46698 149274
rect 46866 149144 47710 149274
rect 47878 149144 48630 149274
rect 48798 149144 49642 149274
rect 49810 149144 50562 149274
rect 50730 149144 51574 149274
rect 51742 149144 52494 149274
rect 52662 149144 53506 149274
rect 53674 149144 54426 149274
rect 54594 149144 55438 149274
rect 55606 149144 56358 149274
rect 56526 149144 57278 149274
rect 57446 149144 58290 149274
rect 58458 149144 59210 149274
rect 59378 149144 60222 149274
rect 60390 149144 61142 149274
rect 61310 149144 62154 149274
rect 62322 149144 63074 149274
rect 63242 149144 64086 149274
rect 64254 149144 65006 149274
rect 65174 149144 66018 149274
rect 66186 149144 66938 149274
rect 67106 149144 67950 149274
rect 68118 149144 68870 149274
rect 69038 149144 69882 149274
rect 70050 149144 70802 149274
rect 70970 149144 71814 149274
rect 71982 149144 72734 149274
rect 72902 149144 73746 149274
rect 73914 149144 74666 149274
rect 74834 149144 75678 149274
rect 75846 149144 76598 149274
rect 76766 149144 77610 149274
rect 77778 149144 78530 149274
rect 78698 149144 79542 149274
rect 79710 149144 80462 149274
rect 80630 149144 81474 149274
rect 81642 149144 82394 149274
rect 82562 149144 83406 149274
rect 83574 149144 84326 149274
rect 84494 149144 85338 149274
rect 85506 149144 86258 149274
rect 86426 149144 87270 149274
rect 87438 149144 88190 149274
rect 88358 149144 89202 149274
rect 89370 149144 90122 149274
rect 90290 149144 91134 149274
rect 91302 149144 92054 149274
rect 92222 149144 93066 149274
rect 93234 149144 93986 149274
rect 94154 149144 94998 149274
rect 95166 149144 95918 149274
rect 96086 149144 96930 149274
rect 97098 149144 97850 149274
rect 98018 149144 98862 149274
rect 99030 149144 99782 149274
rect 99950 149144 100794 149274
rect 100962 149144 101714 149274
rect 101882 149144 102726 149274
rect 102894 149144 103646 149274
rect 103814 149144 104658 149274
rect 104826 149144 105578 149274
rect 105746 149144 106590 149274
rect 106758 149144 107510 149274
rect 107678 149144 108522 149274
rect 108690 149144 109442 149274
rect 480 711 109552 149144
<< metal3 >>
rect 0 149064 800 149184
rect 0 147568 800 147688
rect 0 146072 800 146192
rect 0 144576 800 144696
rect 0 143080 800 143200
rect 0 141584 800 141704
rect 0 140088 800 140208
rect 0 138456 800 138576
rect 0 136960 800 137080
rect 0 135464 800 135584
rect 0 133968 800 134088
rect 0 132472 800 132592
rect 0 130976 800 131096
rect 0 129480 800 129600
rect 0 127848 800 127968
rect 0 126352 800 126472
rect 0 124856 800 124976
rect 0 123360 800 123480
rect 0 121864 800 121984
rect 0 120368 800 120488
rect 0 118872 800 118992
rect 0 117240 800 117360
rect 0 115744 800 115864
rect 0 114248 800 114368
rect 0 112752 800 112872
rect 109200 112344 110000 112464
rect 0 111256 800 111376
rect 0 109760 800 109880
rect 0 108264 800 108384
rect 0 106632 800 106752
rect 0 105136 800 105256
rect 0 103640 800 103760
rect 0 102144 800 102264
rect 0 100648 800 100768
rect 0 99152 800 99272
rect 0 97656 800 97776
rect 0 96024 800 96144
rect 0 94528 800 94648
rect 0 93032 800 93152
rect 0 91536 800 91656
rect 0 90040 800 90160
rect 0 88544 800 88664
rect 0 87048 800 87168
rect 0 85416 800 85536
rect 0 83920 800 84040
rect 0 82424 800 82544
rect 0 80928 800 81048
rect 0 79432 800 79552
rect 0 77936 800 78056
rect 0 76440 800 76560
rect 0 74808 800 74928
rect 0 73312 800 73432
rect 0 71816 800 71936
rect 0 70320 800 70440
rect 0 68824 800 68944
rect 0 67328 800 67448
rect 0 65832 800 65952
rect 0 64200 800 64320
rect 0 62704 800 62824
rect 0 61208 800 61328
rect 0 59712 800 59832
rect 0 58216 800 58336
rect 0 56720 800 56840
rect 0 55224 800 55344
rect 0 53592 800 53712
rect 0 52096 800 52216
rect 0 50600 800 50720
rect 0 49104 800 49224
rect 0 47608 800 47728
rect 0 46112 800 46232
rect 0 44616 800 44736
rect 0 42984 800 43104
rect 0 41488 800 41608
rect 0 39992 800 40112
rect 0 38496 800 38616
rect 109200 37408 110000 37528
rect 0 37000 800 37120
rect 0 35504 800 35624
rect 0 34008 800 34128
rect 0 32376 800 32496
rect 0 30880 800 31000
rect 0 29384 800 29504
rect 0 27888 800 28008
rect 0 26392 800 26512
rect 0 24896 800 25016
rect 0 23400 800 23520
rect 0 21768 800 21888
rect 0 20272 800 20392
rect 0 18776 800 18896
rect 0 17280 800 17400
rect 0 15784 800 15904
rect 0 14288 800 14408
rect 0 12792 800 12912
rect 0 11160 800 11280
rect 0 9664 800 9784
rect 0 8168 800 8288
rect 0 6672 800 6792
rect 0 5176 800 5296
rect 0 3680 800 3800
rect 0 2184 800 2304
rect 0 688 800 808
<< obsm3 >>
rect 880 148984 109200 149157
rect 800 147768 109200 148984
rect 880 147488 109200 147768
rect 800 146272 109200 147488
rect 880 145992 109200 146272
rect 800 144776 109200 145992
rect 880 144496 109200 144776
rect 800 143280 109200 144496
rect 880 143000 109200 143280
rect 800 141784 109200 143000
rect 880 141504 109200 141784
rect 800 140288 109200 141504
rect 880 140008 109200 140288
rect 800 138656 109200 140008
rect 880 138376 109200 138656
rect 800 137160 109200 138376
rect 880 136880 109200 137160
rect 800 135664 109200 136880
rect 880 135384 109200 135664
rect 800 134168 109200 135384
rect 880 133888 109200 134168
rect 800 132672 109200 133888
rect 880 132392 109200 132672
rect 800 131176 109200 132392
rect 880 130896 109200 131176
rect 800 129680 109200 130896
rect 880 129400 109200 129680
rect 800 128048 109200 129400
rect 880 127768 109200 128048
rect 800 126552 109200 127768
rect 880 126272 109200 126552
rect 800 125056 109200 126272
rect 880 124776 109200 125056
rect 800 123560 109200 124776
rect 880 123280 109200 123560
rect 800 122064 109200 123280
rect 880 121784 109200 122064
rect 800 120568 109200 121784
rect 880 120288 109200 120568
rect 800 119072 109200 120288
rect 880 118792 109200 119072
rect 800 117440 109200 118792
rect 880 117160 109200 117440
rect 800 115944 109200 117160
rect 880 115664 109200 115944
rect 800 114448 109200 115664
rect 880 114168 109200 114448
rect 800 112952 109200 114168
rect 880 112672 109200 112952
rect 800 112544 109200 112672
rect 800 112264 109120 112544
rect 800 111456 109200 112264
rect 880 111176 109200 111456
rect 800 109960 109200 111176
rect 880 109680 109200 109960
rect 800 108464 109200 109680
rect 880 108184 109200 108464
rect 800 106832 109200 108184
rect 880 106552 109200 106832
rect 800 105336 109200 106552
rect 880 105056 109200 105336
rect 800 103840 109200 105056
rect 880 103560 109200 103840
rect 800 102344 109200 103560
rect 880 102064 109200 102344
rect 800 100848 109200 102064
rect 880 100568 109200 100848
rect 800 99352 109200 100568
rect 880 99072 109200 99352
rect 800 97856 109200 99072
rect 880 97576 109200 97856
rect 800 96224 109200 97576
rect 880 95944 109200 96224
rect 800 94728 109200 95944
rect 880 94448 109200 94728
rect 800 93232 109200 94448
rect 880 92952 109200 93232
rect 800 91736 109200 92952
rect 880 91456 109200 91736
rect 800 90240 109200 91456
rect 880 89960 109200 90240
rect 800 88744 109200 89960
rect 880 88464 109200 88744
rect 800 87248 109200 88464
rect 880 86968 109200 87248
rect 800 85616 109200 86968
rect 880 85336 109200 85616
rect 800 84120 109200 85336
rect 880 83840 109200 84120
rect 800 82624 109200 83840
rect 880 82344 109200 82624
rect 800 81128 109200 82344
rect 880 80848 109200 81128
rect 800 79632 109200 80848
rect 880 79352 109200 79632
rect 800 78136 109200 79352
rect 880 77856 109200 78136
rect 800 76640 109200 77856
rect 880 76360 109200 76640
rect 800 75008 109200 76360
rect 880 74728 109200 75008
rect 800 73512 109200 74728
rect 880 73232 109200 73512
rect 800 72016 109200 73232
rect 880 71736 109200 72016
rect 800 70520 109200 71736
rect 880 70240 109200 70520
rect 800 69024 109200 70240
rect 880 68744 109200 69024
rect 800 67528 109200 68744
rect 880 67248 109200 67528
rect 800 66032 109200 67248
rect 880 65752 109200 66032
rect 800 64400 109200 65752
rect 880 64120 109200 64400
rect 800 62904 109200 64120
rect 880 62624 109200 62904
rect 800 61408 109200 62624
rect 880 61128 109200 61408
rect 800 59912 109200 61128
rect 880 59632 109200 59912
rect 800 58416 109200 59632
rect 880 58136 109200 58416
rect 800 56920 109200 58136
rect 880 56640 109200 56920
rect 800 55424 109200 56640
rect 880 55144 109200 55424
rect 800 53792 109200 55144
rect 880 53512 109200 53792
rect 800 52296 109200 53512
rect 880 52016 109200 52296
rect 800 50800 109200 52016
rect 880 50520 109200 50800
rect 800 49304 109200 50520
rect 880 49024 109200 49304
rect 800 47808 109200 49024
rect 880 47528 109200 47808
rect 800 46312 109200 47528
rect 880 46032 109200 46312
rect 800 44816 109200 46032
rect 880 44536 109200 44816
rect 800 43184 109200 44536
rect 880 42904 109200 43184
rect 800 41688 109200 42904
rect 880 41408 109200 41688
rect 800 40192 109200 41408
rect 880 39912 109200 40192
rect 800 38696 109200 39912
rect 880 38416 109200 38696
rect 800 37608 109200 38416
rect 800 37328 109120 37608
rect 800 37200 109200 37328
rect 880 36920 109200 37200
rect 800 35704 109200 36920
rect 880 35424 109200 35704
rect 800 34208 109200 35424
rect 880 33928 109200 34208
rect 800 32576 109200 33928
rect 880 32296 109200 32576
rect 800 31080 109200 32296
rect 880 30800 109200 31080
rect 800 29584 109200 30800
rect 880 29304 109200 29584
rect 800 28088 109200 29304
rect 880 27808 109200 28088
rect 800 26592 109200 27808
rect 880 26312 109200 26592
rect 800 25096 109200 26312
rect 880 24816 109200 25096
rect 800 23600 109200 24816
rect 880 23320 109200 23600
rect 800 21968 109200 23320
rect 880 21688 109200 21968
rect 800 20472 109200 21688
rect 880 20192 109200 20472
rect 800 18976 109200 20192
rect 880 18696 109200 18976
rect 800 17480 109200 18696
rect 880 17200 109200 17480
rect 800 15984 109200 17200
rect 880 15704 109200 15984
rect 800 14488 109200 15704
rect 880 14208 109200 14488
rect 800 12992 109200 14208
rect 880 12712 109200 12992
rect 800 11360 109200 12712
rect 880 11080 109200 11360
rect 800 9864 109200 11080
rect 880 9584 109200 9864
rect 800 8368 109200 9584
rect 880 8088 109200 8368
rect 800 6872 109200 8088
rect 880 6592 109200 6872
rect 800 5376 109200 6592
rect 880 5096 109200 5376
rect 800 3880 109200 5096
rect 880 3600 109200 3880
rect 800 2384 109200 3600
rect 880 2104 109200 2384
rect 800 888 109200 2104
rect 880 715 109200 888
<< metal4 >>
rect 4208 2128 4528 147472
rect 19568 2128 19888 147472
rect 34928 2128 35248 147472
rect 50288 2128 50608 147472
rect 65648 2128 65968 147472
rect 81008 2128 81328 147472
rect 96368 2128 96688 147472
<< obsm4 >>
rect 1715 3979 4128 147117
rect 4608 3979 19488 147117
rect 19968 3979 34848 147117
rect 35328 3979 50208 147117
rect 50688 3979 65568 147117
rect 66048 3979 80928 147117
rect 81408 3979 96288 147117
rect 96768 3979 105925 147117
<< labels >>
rlabel metal2 s 478 149200 534 150000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 29366 149200 29422 150000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 32310 149200 32366 150000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 35162 149200 35218 150000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 38106 149200 38162 150000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 40958 149200 41014 150000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 43902 149200 43958 150000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 46754 149200 46810 150000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 49698 149200 49754 150000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 52550 149200 52606 150000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 55494 149200 55550 150000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3330 149200 3386 150000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 58346 149200 58402 150000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 61198 149200 61254 150000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 64142 149200 64198 150000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 66994 149200 67050 150000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 69938 149200 69994 150000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 72790 149200 72846 150000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 75734 149200 75790 150000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 78586 149200 78642 150000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 81530 149200 81586 150000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 84382 149200 84438 150000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6182 149200 6238 150000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 87326 149200 87382 150000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 90178 149200 90234 150000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 93122 149200 93178 150000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 95974 149200 96030 150000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 98918 149200 98974 150000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 101770 149200 101826 150000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 104714 149200 104770 150000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 107566 149200 107622 150000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9126 149200 9182 150000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 11978 149200 12034 150000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 14922 149200 14978 150000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 17774 149200 17830 150000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 20718 149200 20774 150000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 23570 149200 23626 150000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 26514 149200 26570 150000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1398 149200 1454 150000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 30378 149200 30434 150000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 33230 149200 33286 150000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 36174 149200 36230 150000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 39026 149200 39082 150000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 41970 149200 42026 150000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 44822 149200 44878 150000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 47766 149200 47822 150000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 50618 149200 50674 150000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 53562 149200 53618 150000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 56414 149200 56470 150000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 4250 149200 4306 150000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 59266 149200 59322 150000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 62210 149200 62266 150000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 65062 149200 65118 150000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 68006 149200 68062 150000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 70858 149200 70914 150000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 73802 149200 73858 150000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 76654 149200 76710 150000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 79598 149200 79654 150000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 82450 149200 82506 150000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 85394 149200 85450 150000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 7194 149200 7250 150000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 88246 149200 88302 150000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 91190 149200 91246 150000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 94042 149200 94098 150000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 96986 149200 97042 150000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 99838 149200 99894 150000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 102782 149200 102838 150000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 105634 149200 105690 150000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 108578 149200 108634 150000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 10046 149200 10102 150000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 12990 149200 13046 150000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 15842 149200 15898 150000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 18786 149200 18842 150000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 21638 149200 21694 150000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 24582 149200 24638 150000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 27434 149200 27490 150000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2318 149200 2374 150000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 31298 149200 31354 150000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 34242 149200 34298 150000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 37094 149200 37150 150000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 40038 149200 40094 150000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 42890 149200 42946 150000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 45834 149200 45890 150000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 48686 149200 48742 150000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 51630 149200 51686 150000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 54482 149200 54538 150000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 57334 149200 57390 150000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 5262 149200 5318 150000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 60278 149200 60334 150000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 63130 149200 63186 150000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 66074 149200 66130 150000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 68926 149200 68982 150000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 71870 149200 71926 150000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 74722 149200 74778 150000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 77666 149200 77722 150000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 80518 149200 80574 150000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 83462 149200 83518 150000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 86314 149200 86370 150000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 8114 149200 8170 150000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 89258 149200 89314 150000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 92110 149200 92166 150000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 95054 149200 95110 150000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 97906 149200 97962 150000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 100850 149200 100906 150000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 103702 149200 103758 150000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 106646 149200 106702 150000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 109498 149200 109554 150000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 11058 149200 11114 150000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 13910 149200 13966 150000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 16854 149200 16910 150000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 19706 149200 19762 150000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 22650 149200 22706 150000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 25502 149200 25558 150000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 28446 149200 28502 150000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 109200 37408 110000 37528 6 la_blink[0]
port 115 nsew signal output
rlabel metal3 s 109200 112344 110000 112464 6 la_blink[1]
port 116 nsew signal output
rlabel metal4 s 4208 2128 4528 147472 6 vccd1
port 117 nsew power input
rlabel metal4 s 34928 2128 35248 147472 6 vccd1
port 117 nsew power input
rlabel metal4 s 65648 2128 65968 147472 6 vccd1
port 117 nsew power input
rlabel metal4 s 96368 2128 96688 147472 6 vccd1
port 117 nsew power input
rlabel metal4 s 19568 2128 19888 147472 6 vssd1
port 118 nsew ground input
rlabel metal4 s 50288 2128 50608 147472 6 vssd1
port 118 nsew ground input
rlabel metal4 s 81008 2128 81328 147472 6 vssd1
port 118 nsew ground input
rlabel metal3 s 0 688 800 808 6 wb_ack_o
port 119 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 wb_adr_i[0]
port 120 nsew signal input
rlabel metal3 s 0 62704 800 62824 6 wb_adr_i[10]
port 121 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 wb_adr_i[11]
port 122 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 wb_adr_i[12]
port 123 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 wb_adr_i[13]
port 124 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 wb_adr_i[14]
port 125 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 wb_adr_i[15]
port 126 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 wb_adr_i[16]
port 127 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 wb_adr_i[17]
port 128 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 wb_adr_i[18]
port 129 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 wb_adr_i[19]
port 130 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 wb_adr_i[1]
port 131 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 wb_adr_i[20]
port 132 nsew signal input
rlabel metal3 s 0 112752 800 112872 6 wb_adr_i[21]
port 133 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 wb_adr_i[22]
port 134 nsew signal input
rlabel metal3 s 0 121864 800 121984 6 wb_adr_i[23]
port 135 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 wb_adr_i[2]
port 136 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 wb_adr_i[3]
port 137 nsew signal input
rlabel metal3 s 0 35504 800 35624 6 wb_adr_i[4]
port 138 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 wb_adr_i[5]
port 139 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 wb_adr_i[6]
port 140 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 wb_adr_i[7]
port 141 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 wb_adr_i[8]
port 142 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 wb_adr_i[9]
port 143 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wb_clk_i
port 144 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 wb_cyc_i
port 145 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 wb_data_i[0]
port 146 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 wb_data_i[10]
port 147 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 wb_data_i[11]
port 148 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 wb_data_i[12]
port 149 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 wb_data_i[13]
port 150 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 wb_data_i[14]
port 151 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 wb_data_i[15]
port 152 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 wb_data_i[16]
port 153 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 wb_data_i[17]
port 154 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 wb_data_i[18]
port 155 nsew signal input
rlabel metal3 s 0 105136 800 105256 6 wb_data_i[19]
port 156 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 wb_data_i[1]
port 157 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 wb_data_i[20]
port 158 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 wb_data_i[21]
port 159 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 wb_data_i[22]
port 160 nsew signal input
rlabel metal3 s 0 123360 800 123480 6 wb_data_i[23]
port 161 nsew signal input
rlabel metal3 s 0 126352 800 126472 6 wb_data_i[24]
port 162 nsew signal input
rlabel metal3 s 0 129480 800 129600 6 wb_data_i[25]
port 163 nsew signal input
rlabel metal3 s 0 132472 800 132592 6 wb_data_i[26]
port 164 nsew signal input
rlabel metal3 s 0 135464 800 135584 6 wb_data_i[27]
port 165 nsew signal input
rlabel metal3 s 0 138456 800 138576 6 wb_data_i[28]
port 166 nsew signal input
rlabel metal3 s 0 141584 800 141704 6 wb_data_i[29]
port 167 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 wb_data_i[2]
port 168 nsew signal input
rlabel metal3 s 0 144576 800 144696 6 wb_data_i[30]
port 169 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 wb_data_i[31]
port 170 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 wb_data_i[3]
port 171 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 wb_data_i[4]
port 172 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 wb_data_i[5]
port 173 nsew signal input
rlabel metal3 s 0 46112 800 46232 6 wb_data_i[6]
port 174 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 wb_data_i[7]
port 175 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 wb_data_i[8]
port 176 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 wb_data_i[9]
port 177 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 wb_data_o[0]
port 178 nsew signal output
rlabel metal3 s 0 65832 800 65952 6 wb_data_o[10]
port 179 nsew signal output
rlabel metal3 s 0 70320 800 70440 6 wb_data_o[11]
port 180 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 wb_data_o[12]
port 181 nsew signal output
rlabel metal3 s 0 79432 800 79552 6 wb_data_o[13]
port 182 nsew signal output
rlabel metal3 s 0 83920 800 84040 6 wb_data_o[14]
port 183 nsew signal output
rlabel metal3 s 0 88544 800 88664 6 wb_data_o[15]
port 184 nsew signal output
rlabel metal3 s 0 93032 800 93152 6 wb_data_o[16]
port 185 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 wb_data_o[17]
port 186 nsew signal output
rlabel metal3 s 0 102144 800 102264 6 wb_data_o[18]
port 187 nsew signal output
rlabel metal3 s 0 106632 800 106752 6 wb_data_o[19]
port 188 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 wb_data_o[1]
port 189 nsew signal output
rlabel metal3 s 0 111256 800 111376 6 wb_data_o[20]
port 190 nsew signal output
rlabel metal3 s 0 115744 800 115864 6 wb_data_o[21]
port 191 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 wb_data_o[22]
port 192 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 wb_data_o[23]
port 193 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 wb_data_o[24]
port 194 nsew signal output
rlabel metal3 s 0 130976 800 131096 6 wb_data_o[25]
port 195 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 wb_data_o[26]
port 196 nsew signal output
rlabel metal3 s 0 136960 800 137080 6 wb_data_o[27]
port 197 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 wb_data_o[28]
port 198 nsew signal output
rlabel metal3 s 0 143080 800 143200 6 wb_data_o[29]
port 199 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 wb_data_o[2]
port 200 nsew signal output
rlabel metal3 s 0 146072 800 146192 6 wb_data_o[30]
port 201 nsew signal output
rlabel metal3 s 0 149064 800 149184 6 wb_data_o[31]
port 202 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 wb_data_o[3]
port 203 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 wb_data_o[4]
port 204 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 wb_data_o[5]
port 205 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 wb_data_o[6]
port 206 nsew signal output
rlabel metal3 s 0 52096 800 52216 6 wb_data_o[7]
port 207 nsew signal output
rlabel metal3 s 0 56720 800 56840 6 wb_data_o[8]
port 208 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 wb_data_o[9]
port 209 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 wb_rst_i
port 210 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wb_sel_i[0]
port 211 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 wb_sel_i[1]
port 212 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 wb_sel_i[2]
port 213 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 wb_sel_i[3]
port 214 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 wb_stall_o
port 215 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 wb_stb_i
port 216 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 wb_we_i
port 217 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 110000 150000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 45637670
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripherals_Flat/runs/Peripherals_Flat/results/finishing/Peripherals.magic.gds
string GDS_START 1229070
<< end >>

